En hjälp ville lägga om ett foto journalist frågade den retoriska frågan:Om du befunnit dig i en situation där du kan antingen sparaen drunknande, eller du kan ta en Pulitzer prisvinnandefotografi av honom drunkning, vilken slutarhastighet och inställning skulle du använda?
		-- Paul Harvey

%
En höna Ruvande KattungarEn vän berättar att han såg i Novato ranch, Marin County,några dagar sedan, en höna faktiskt ruvande och annat hand om trekattungar! The gentleman på vars lokaler denna märkliga händelse transpiringsäger hönan antog ungarna när de var men några dagar gammal, och attHon har ägnat dem sin odelade vård för flera veckor tidigare. De ungakattdjur är nu av respektabel storlek, men de ändå följa hönan påhennes cluckings och regelbundet grubblat på natten under sina vingar.
		-- Sacramento Daily Union, July 2, 1861

%
En journalist, glada över sin middag, frågade kocken för receptet.Svarade kocken, "Vi har samma politik som ni journalister, vialdrig avslöja vår sås. "
		-- Sacramento Daily Union, July 2, 1861

%
En mexikansk tidning rapporterar att uttråkade Royal Air Force piloter stationepå Falklandsöarna har utarbetat vad de anser en fantastisk nyspel. Notera att de lokala pingviner är fascinerad av flygplan, denpiloter söker en strand där fåglarna samlas och flyga långsamtlängs den i vattnet. Kanske tiotusen pingviner vända derashuvuden unisont tittar på planen går, och när piloterna vändarunt och flyga tillbaka, fåglarna vända huvudet i motsattriktning, som åskådare vid en slow-motion tennismatch. Sedanpappersrapporter "Piloterna flyger ut till havs och direkt till pingvinenkoloni och flyga den. Heads gå upp, upp, upp, och tio tusen pingvinerfalla försiktigt på ryggen.
		-- Audobon Society Magazine

%
Ett nytt sätt att ta pillerEn läkare en natt i Wisconsin störs av en inbrottstjuv, ochhar ingen boll eller skott för hans pistol, ljudlöst laddade vapnet medsmå, hårda piller och gav inkräktaren ett "recept", som han tyckerkommer att gå långt mot härdning rascalen av en mycket dålig krämpa.
		-- Nevada Morning Transcript, January 30, 1861

%
En tidning är en cirkulerande bibliotek med högt blodtryck.
		-- Arthure "Bugs" Baer

%
En framstående program på en storvilts safari i Afrika, fördes till envattenhål där kunde observeras livet i djungeln. När hantittade ner från sitt träd plattform och beskrev scenen i sinbandspelare, såg han två gnuer betar fredligt. Så upptagen varde att de åsidosatt en metod med en stolthet av lejon leddemed två magnifika exemplar, uppenbarligen ledarna. Lejon laddade,dödade gnuer, och släpade dem in i buskarna där deras festandekunde inte ses. En liten stund senare de två kungarna i djungelnuppstått och radioman inspelad på hans band: "Ja, det är i slutet avden gnus och här, återigen, är de huvud lejon. "
		-- Arthure "Bugs" Baer

%
"En tvättbjörn trassla med en 23.000 volt nätet idag. Resultaten blackoutut 1400 bostäder och, naturligtvis, en tvättbjörn. "
		-- Steel City News

%
En ung flicka en gång begått självmord eftersom hennes mamma vägrade henne en nyhätta. Coroner dom: "Död från överdriven spunk."
		-- Sacramento Daily Union, September 13, 1860

%
Annonser innehåller de enda sanningar för att kunna åberopas i en tidning.
		-- Thomas Jefferson

%
Efter två eller tre veckor av denna galenskap, börjar du känna ett medmannen som sade, "Inga nyheter är goda nyheter." I tjugoåtta papper, endastden mest sällsynta typen av lycka kommer att dyka upp mer än två eller tre artiklarnågot intresse ... men även då de ränteposter vanligen begravda djuptrunt punkt 16 på hoppet (eller "Forts. på ...") sida ...Posten kommer att ha en historia om Muskie ett tal i Iowa. DeStar kommer att säga samma sak, och Journal säger ingenting alls.Men tiderna kan ha tillräckligt med utrymme på hoppet för att inkludera en radeller så som säger något i stil med: "När han avslutade sitt tal, Muskiebrast i gråt och grep hans kampanjledare vid sidan av halsen.De brottats kort, men kampen sparkades sönder av en orientaliskkvinna som verkade ha kontroll. "Nu det är bra journalistik. Helt mål; mycket aktiv och raktill poängen.
		-- Hunter S. Thompson, "Fear and Loathing '72"

%
Alla tidningen ledarskribenter någonsin göra är att komma ned från bergen efterstriden är över och skjuta den sårade.
		-- Hunter S. Thompson, "Fear and Loathing '72"

%
En redaktör är en som skiljer agnarna från vetet och skriver vetet.
		-- Adlai Stevenson

%
"... Och kom ihåg: om du inte gillar nyheter, gå ut och göra en del avdin egen."
		-- "Scoop" Nisker, KFOG radio reporter Preposterous Words

%
Och det är så det är ...
		-- Walter Cronkite

%
Jorden förstörd av Solar Flare - filmklipp på elva.
		-- Walter Cronkite

%
Varje journalist har en roman i sig, vilket är en utmärkt plats för det.
		-- Walter Cronkite

%
Allt du läser i tidningar är helt sant, med undantag för detsällsynt berättelse som du råkar ha förstahandsinformation.
		-- Erwin Knoll

%
BLIXT!Intelligens av mänskligheten minskar.Detaljer på ... eh, när den lilla handen är på ....
		-- Erwin Knoll

%
... Hade detta varit en verklig nödsituation, vi skulle ha flytt i skräck,och du inte skulle ha underrättats.
		-- Erwin Knoll

%
Jag vet bara vad jag läst i tidningarna.
		-- Will Rogers

%
Jag läser tidningen glupskt. Det är min en form av kontinuerlig fiction.
		-- Aneurin Bevan

%
Jag ser verkligen med medömkan över den stora kroppen av mina landsmänsom läser tidningar, leva och dö i tron ​​att de har käntnågot av vad som har passerat på sin tid.
		-- H. Truman

%
Om jag skulle gå på vatten, skulle pressen säga att jag bara gör deteftersom jag kan inte simma.
		-- Bob Stanfield

%
Om du tappar humöret på en tidningskåsör, kommer han bli rik,eller känd eller båda.
		-- Bob Stanfield

%
I ett medium i vilket en nyhets Piece tar en minut och en "djupgående"Piece tar två minuter, kommer Simple driva ut komplexet.
		-- Frank Mankiewicz

%
Är det inte tänkbart för er att en intelligent person kan hysatvå motsatta idéer i hans sinne?
		-- Adlai Stevenson, to reporters

%
Dess brister Trots det finns mycket att säga till förmån för journalistiki det genom att ge oss yttrandet från outbildade, det håller oss i kontakt medokunnighet i samhället.
		-- Oscar Wilde

%
Journalistik är litteratur bråttom.
		-- Matthew Arnold

%
Journalistik kommer att döda dig, men det kommer att hålla dig vid liv när du ändå håller på.
		-- Matthew Arnold

%
De flesta berg journalistik är människor som inte kan skriva intervjua människor somkan inte tala för människor som inte kan läsa.
		-- Frank Zappa

%
Min far var en gudfruktig man, men han missade aldrig en kopia avNew York Times, heller.
		-- E. B. White

%
förolämpa aldrig människor med stil när du kan förolämpa dem med ämnet.
		-- Sam Brown, "The Washington Post", January 26, 1977

%
   *** Inforuta ***Ryska stridsvagnar steamrolling genom New Jersey !!!! Detaljer på elva!
		-- Sam Brown, "The Washington Post", January 26, 1977

%
"Ingen självaktning fisk vill vara insvept i den typen av papper."övertas av Rupert Murdoch
		-- Mike Royko on the Chicago Sun-Times after it was

%
Av vad du ser i böcker, tror 75%. Tidningar, tror 50%. ochTV-nyheter, tror 25% - göra det 5% om ankare bär en kavaj.
		-- Mike Royko on the Chicago Sun-Times after it was

%
Än en gång UppifrånKorrigering meddelande i Miami Herald: "I söndags The Herald felaktigtrapporterade den ursprungliga Dolphin Johnny Holmes hade varit en försäkring försäljarei Raleigh, North Carolina, att han hade vunnit New York lotteri 1982 ochförlorade pengar i ett land svindel, att han hade åtalats för fordonstrafikmord, men frikändes eftersom hans mamma sa att hon körde bilen, och attHan uppgav att det roligaste han någonsin såg var Flipper sprutande vatten påGeorge Wilson. Var och en av dessa poster var felaktiga material som publicerasoavsiktligt. Han var inte en försäkring försäljare i Raleigh, inte vinnalotteri, var varken han eller hans mor laddade eller på något sätt har medvehicular homicide, och han gjorde ingen kommentar om Flipper eller George Wilson.Herald beklagar felen. "
		-- "The Progressive", March, 1987

%
Ett av tecknen på Napoleons storhet är det faktum att han en gång hade enutgivare skott.
		-- Siegfried Unseld

%
Människor som är roliga och smarta och retur telefonsamtal får mycket bättretryck än människor som är bara roligt och smart.
		-- Howard Simons, "The Washington Post"

%
Fotografera en vulkan är bara om de mest eländiga sak du kan göra.[Vem har uppenbarligen aldrig försökt att använda en PDP-10. Ed.]
		-- Robert B. Goodman

%
Reportrar som Bill Greider från Washington Post och HimNaughton i New York Times, till exempel, var tvungen att lämna långa, detaljerade,och relativt komplexa berättelser varje dag - medan min egen deadline föllvarannan vecka - men ingen av dem någonsin verkade bråttom omfå jobbet gjort, och från tid till tid de skulle försöka tröstamig om den fruktansvärda trycket jag alltid tycktes vara arbetande under.Alla $ 100 en timme psykiater kan nog förklara detta problemtill mig, i tretton eller fjorton sessioner, men jag har inte tid för det.Ingen tvekan om det har något att göra med en djupt rotad personlighet defekt, ellerkanske en knut i vilken blodkärlet leder till tallkottkörteln ... PåDäremot kan det vara något så enkelt och i princip perversa somoavsett instinkt är det som orsakar en jackrabbit att vänta tills den sistaeventuella andra att dart tvärs över vägen framför bilen fortkörning.
		-- Hunter S. Thompson, "Fear and Loathing on the Campaign Trail"

%
Annonsen är den mest sannfärdiga delen i en tidning.
		-- Thomas Jefferson

%
American Dental Association meddelade idag att de flesta plack tenderarbildas på tänderna runt 4:00 på eftermiddagen.Film på 11:00.
		-- Thomas Jefferson

%
Den viktigaste tjänsten utförs av pressen är att utbildamänniskor att närma trycksaker med misstro.
		-- Thomas Jefferson

%
"The New York Times läses av människor som driver landet. DenWashington Post läses av människor som tror att de kör landet. DeNational Enquirer läses av människor som tror att Elvis lever och körlandet ..."
		-- Robert J Woodhead

%
De enda egenskaper för verklig framgång i journalistik är ratlike list, enrimligt sätt och en liten litterär förmåga. Förmågan att stjälaandras idéer och fraser ... är också ovärderligt.
		-- Nicolas Tomalin, "Stop the Press, I Want to Get On"

%
Världen är verkligen inte något värre. Det är bara det att nyhetsbevakningenär så mycket bättre.
		-- Nicolas Tomalin, "Stop the Press, I Want to Get On"

%
"Då du erkänner som bekräftar inte förneka du någonsin sagt det?""NEJ! ... Jag menar Ja! VAD?""Jag ska sätta` kanske. "
		-- Bloom County

%
Detta är ett test av den akuta sändningssystem. Hade det funnits enverklig nödsituation, då skulle du inte längre här.
		-- Bloom County

%
Detta är ett test av Emergency Broadcast System. Om detta hade varit enverklig nödsituation, tror du verkligen att vi skulle stanna kvar för att berätta?
		-- Bloom County

%
Detta liv är ett test. Det är bara ett test. Hade detta varit ett verkliga livet, duskulle ha fått ytterligare instruktioner om vad man ska göra och vart den ska gå.
		-- Bloom County

%
Varning: Lyssna på WXRT på första april rekommenderas inte förde som är något förvirrade de första timmarna efter uppvaknandet.
		-- Chicago Reader 4/22/83

%
Du vet den stora sak om TV? Om något viktigt händernågonstans alls i världen, oavsett vilken tid på dagen eller natten,Du kan alltid byta kanal.
		-- Jim Ignatowski

%
