En baby är en matsmältningskanalen med hög röst i ena änden och ingenansvar i den andra.
		-- George Bernard Shaw

%
En baby är Guds yttrande att världen bör gå på.
		-- Carl Sandburg

%
Ett barn av fem kunde förstå detta! Hämta mig ett barn av fem.
		-- Carl Sandburg

%
En kid'll äta mitt i en Oreo, så småningom.
		-- Carl Sandburg

%
Ett litet barn gick upp till Santa och frågade honom: "Santa, du vet när jag är dåligeller hur? "Och Santa säger:" Ja, det gör jag. "Den lilla ungen frågar då:" Och duvet när jag sover? "Till vilken Santa svarar:" Varje minut. "Sålitet barn säger då, "Ja, om du vet när jag är dålig och när jag är bra,hur kommer du inte vet vad jag vill ha i julklapp? "
		-- Carl Sandburg

%
Ett ungt gift par hade sitt första barn. Deras ursprungliga stolthetoch glädje vände sig långsamt till oro men för efter ett par år debarn hade aldrig yttrat någon form av tal. De anlitade bästa talterapeuter, läkare, psykiatriker, alla förgäves. Barnet helt enkelt vägratatt tala. En morgon när barnet var fem, medan mannen lästepapperet, och hustrun var utfodring hunden, ser den lilla ungen upp frånsin skål och sa, "Min spannmål kallt."Paret är chockad. Mannen, i tårar, konfronterar sin son. "Son,efter alla dessa år, varför har du väntat så länge med att säga något? ".Rycker ungen, "Allt har varit okej 'til nu".
		-- Carl Sandburg

%
Om det enda vi har kvar som faktiskt diskriminerar till förmån förde vanligt folk är storken.
		-- Carl Sandburg

%
Adam och Eva hade många fördelar, men den huvudsakliga var att de flyddetandsprickning.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Adopterade barn är en sådan smärta - man måste lära dem att se ut som du ...
		-- Gilda Radner

%
Efter att ha sett en mycket attraktiv mamma ward patientenuppriktigt tumme sig igenom en telefonkatalog för fleraminuter, ett sjukhus ordnad slutligen frågade om han kunde vara till någon hjälp."Nej tack", log den unga modern, "Jag är bara ute efter ennamn för mitt barn. ""Men sjukhuset levererar en särskild broschyr som listar hundratalsförsta namn och deras betydelser ", sade ordnad."Det kommer inte att hjälpa", sade kvinnan, "mitt barn har redan ett förnamn."
		-- Gilda Radner

%
Och han klättrade med lad upp Eiffelberg Tower. "Detta", ropade borgmästaren,"Är din stad mörkaste timme! Tiden för alla Whos som har blod som är röttatt komma till hjälp av deras land! ", sade han." Vi har att göra ljud istörre mängder! Så, öppna munnen, gosse! För varje röst räknas! "Så hantalade som han klättrade. När de kom till toppen, pojken harklade sig ochHan ropade, "YOPP!"Och att Yopp ... Att en sista liten, extra Yopp placera den över!Slutligen, äntligen! Från fläck på den klöver deras röster hördes!De ringde ut klart och rent. Och de elefant log. "Ser du vadJag menar? "De har visat att de är personer, oavsett hur liten. Och derashela världen räddades av den minsta av alla! ""Hur sant! Ja, hur sant", sade den stora känguru. "Och från och med nupå, vet du vad jag planerar att göra? Från och med nu kommer jag att skyddadem med dig! "Och den unge känguru i sin påse sade," me too! Frånsolen på sommaren. Från regn när det är höst-ish, jag kommer att skyddadem. Oavsett hur små-ish! "
		-- Dr. Seuss "Horton Hears a Who"

%
Alla far som tror att han är alla viktiga bör påminna sig om att dettalands hedrar fäder endast en dag om året medan pickles få en hel vecka.
		-- Dr. Seuss "Horton Hears a Who"

%
Alla som använder frasen "enkelt som att ta godis från ett barn" har aldrigförsökte ta godis från ett barn.
		-- Robin Hood

%
Är du förälder? Har du ibland själv osäker på vadsäger i dessa besvärliga situationer? Oroa dig inte mer ...Är du säker på att berätta att du sanningen? Tänk hårt.Gör det dig glad att veta att du skickar mig till en tidig död?Om alla dina vänner hoppade av klippan, skulle du hoppa också?Känner du dig illa? Hur tror du jag känner?Är du inte skämmas?Vet du inte bättre?Hur kan du vara så dum?Om det är det värsta smärta du någonsin kommer att känna, bör du vara tacksamma.Du kan inte lura mig. Jag vet vad du tänker.Om du inte kan säga något trevligt, säger ingenting alls.
		-- Robin Hood

%
Är du förälder? Har du ibland själv osäker på vadsäger i dessa besvärliga situationer? Oroa dig inte mer ...Gör som jag säger, inte som jag gör.Gör mig en tjänst och inte berätta om det. Jag vill inte veta.Vad gjorde du * här * tid?Om det inte smaka illa, skulle det inte vara bra för dig.När jag var i din ålder ...Jag kommer inte älska dig om du fortsätter att göra det.Tänk på alla svältande barn i Indien.Om det finns en sak som jag hatar, det är en lögnare.	Jag ska döda dig.Way to go, klumpig.Om du inte gillar det, kan du bunta det.
		-- Robin Hood

%
Är du förälder? Har du ibland själv osäker på vadsäger i dessa besvärliga situationer? Oroa dig inte mer ...Gå bort. Du bry mig.	Varför? Eftersom livet är orättvist.Det är en fin teckning. Vad är det?Barn ska ses men inte höras.Du kommer att vara död mig.Du kommer att förstå när du blir äldre.	Därför att.Torka den leende utanför ditt ansikte.Jag tror inte du.Hur många gånger har jag sagt till dig att vara försiktig?	Bara för att.
		-- Robin Hood

%
Är du förälder? Har du ibland själv osäker på vadsäger i dessa besvärliga situationer? Oroa dig inte mer ...Bra barn alltid lyda.Sluta agerar så barnslig.Pojkar gråter inte.Om du fortsätta att göra ansikten, en dag det kommer att frysa på det sättet.Varför har du att veta så mycket?Detta skadar mig mer än det skadar dig.	Varför? Eftersom jag är större än du.Tja, har du förstört allt. Nu är du nöjd?Åh, växa upp.Jag bara gör detta eftersom jag älskar dig.
		-- Robin Hood

%
Är du förälder? Har du ibland själv osäker på vadsäger i dessa besvärliga situationer? Oroa dig inte mer ...När kommer ni att växa upp?Jag bara gör det för ditt eget bästa.	Varför gråter du? Sluta gråta, eller jag ska ge dig något attgråta över.Vad är det med dig?En dag du kommer att tacka mig för detta.Du skulle tappa huvudet om det inte var fästa.Inte du har någon mening alls?Om du håller suga tummen, kommer det att falla bort.	Varför? För att jag sa det.Jag hoppas att ni har ett barn precis som dig själv.
		-- Robin Hood

%
Är du förälder? Har du ibland själv osäker på vadsäger i dessa besvärliga situationer? Oroa dig inte mer ...Du skulle inte förstå.Du frågar för många frågor.För att vara en man, måste du lära dig att följa order.Det är för mig att veta och dig att ta reda på.Låt inte dessa mobbare skjuta dig runt. Gå in där och hållaupp för dig själv.Du agerar för stort för dina britches.Tja, bröt du det. Nu är du nöjd?Vänta tills din far kommer hem.Uttråkad? Om du är uttråkad, har jag fått några sysslor för dig.Shape upp eller skicka ut.
		-- Robin Hood

%
Artikel tredje:Om ett brott av njurarna har ägt rum, den tilltalade börha rätt till en snabb blöjbyte. Offentliga tillkännagivanden ochguidade turer i den tidigare nämnda är inte nödvändigt.Artikel fjärde:Beslutet att äta ansträngda lamm eller inte bör vara med "feedee"och inte "feeder". Blåsa ansträngda lamm i mataren sansikte bör accepteras som ett yttrande, inte som en krigsförklaring.Artikel femte:Spädbarn bör njuta av friheten att artikulera, vare sig det är i kyrkan,en offentlig mötesplats under en film, eller efter timmar närljuset är släckt. De har ännu inte lärt sig att glädje och skratt harpågå under en livstid och måste bevaras.
		-- Erma Bombeck, "A Baby's Bill of Rights"

%
Slå din son varje dag; du kanske inte vet varför, men han kommer.
		-- Erma Bombeck, "A Baby's Bill of Rights"

%
Eftersom vi inte tänker på kommande generationer, kommer de aldrig att glömma oss.
		-- Henrik Tikkanen

%
Billy: Mamma, vet du att vasen du sa avkunnades frångeneration till generation?Mamma: Ja?Billy: Tja, denna generation tappade den.
		-- Henrik Tikkanen

%
Amning bör inte försökas av fäder med håriga bröst,eftersom de kan göra barnet nysning och ge den vind.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Fånga hans barn med sina händer i det nya, fortfarande är våt, uteplats,fadern förlorade dem. Hans fru frågade: "Har du inte älskar dina barn?""I det abstrakta, ja, men inte i betongen."
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Catproof är en oxymoron, barn nästan så.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Barn är som katter, kan de säga när du inte gillar dem. det ärnär de kommer över och bryter kroppen utrymme.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Barn är naturliga härmar som fungerar som sina föräldrar trots allaförsök att lära dem gott uppförande.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Barn är oförutsägbara. Man vet aldrig vad inkonsekvens de ärkommer att fånga dig i nästa.
		-- Franklin P. Jones

%
Barn börjar genom att älska sina föräldrar. Efter en tid som de bedömer dem.Sällan, om någonsin, de förlåter dem.
		-- Oscar Wilde

%
Barn sällan felciterar dig. Faktum är att de vanligtvis upprepa ord förord vad du inte borde ha sagt.
		-- Oscar Wilde

%
Barns talang att uthärda härrör från deras okunnighet om alternativ.
		-- Maya Angelou, "I Know Why the Caged Bird Sings"

%
Städning ditt hus medan barnen växer fortfarande är som skottapromenad innan det slutar snöa.Det finns ingen anledning att göra något hushållsarbete alls. Efter de första fyra årensmutsen inte bli värre.
		-- Quentin Crisp

%
Vanföreställningar är ofta funktionella. En mors åsikter om hennes barnsskönhet, intelligens, godhet, et cetera ad nauseam, hålla henne från drunkningdem vid födseln.
		-- Robert Heinlein

%
Inte handikapp dina barn genom att göra deras liv enkelt.
		-- Robert Heinlein

%
Fertilitet är ärftlig. Om dina föräldrar inte har några barn,inte heller kommer du.
		-- Robert Heinlein

%
För vuxenutbildningen inget slår barn.
		-- Robert Heinlein

%
För barn med kort uppmärksamhet spänner: bumeranger som inte kommer tillbaka.
		-- Robert Heinlein

%
FORTUNE MINNS DE STORA FOSTRAR: # 5"Och, och, och, och, men, men, men, men!"
		-- Mrs. Janice Markowsky, April 8, 1965

%
FORTUNE MINNS DE STORA FOSTRAR: # 6"Johnny, om du faller och bryter benet, inte komma springande till mig!"
		-- Mrs. Emily Barstow, June 16, 1954

%
Hämnas! Leva länge nog för att vara ett problem för dina barn!
		-- Mrs. Emily Barstow, June 16, 1954

%
Detta är lätt. Du behöver aldrig räkna ut vad du får för barn,eftersom de kommer att berätta exakt vad de vill. De tillbringar månader ochmånader forskar dessa typer av saker genom att titta på lördag morgontecknad visa annonser. Se till att du får dina barn exakt vadde frågar efter, även om du ogillar deras val. Om ditt barn tänkerhan vill Mord Bob, dockan med ansiktet du kan rippa Rätt off, skulle dubättre få det. Du kan vara orolig att det kan bidra till att uppmuntra dinbarns asociala tendenser, men tro mig, du har inte sett antisocialtendenser tills du har sett ett barn som är övertygad om att han eller hon intefå rätt gåva.
		-- Dave Barry, "Christmas Shopping: A Survivor's Guide"

%
Ge en liten pojke en hammare och han kommer att tycka att allt han stöterbehöver bultande.
		-- Dave Barry, "Christmas Shopping: A Survivor's Guide"

%
Ge ditt barn mentala blockeringar för jul.
		-- Dave Barry, "Christmas Shopping: A Survivor's Guide"

%
Att ha barn är som att ha en bowlingbana installerad i din hjärna.
		-- Martin Mull

%
Hur skarpare än en orm tand är en syster "Ser ni?"
		-- Linus Van Pelt

%
"Humpf!" Humpfed en röst! "För nästan två dagar du har flöda och insisterade påchatta med personer som aldrig existerat. Sådana transporter-on i vår fredligadjungel! Vi har fått nog av er böla bungle! Och jag är här för attstat "brast den stora känguru," Att din fåniga nonsens spelet handlarGenom "Och den unge känguru i sin påse sade," Jag också! ""Med hjälp av Wickersham Brothers och dussintals WickershamMorbröder och Wickersham kusiner och Wickersham svärföräldrar, vars hjälp jag har engagerad,Du kommer att vara avgränsades! Och du kommer att bli bur! Och som för din dammspeck ... Hah! Att vi ska koka i en varm ångande kittel med Beezle-mutter olja! "
		-- Dr. Seuss "Horton Hears a Who"

%
Jag satsar när Neanderthal barn skulle göra en snögubbe, någon skulle alltidsluta säga, "Glöm inte de tjocka tunga ögonbrynen." Då skulle de fågenerad eftersom de ihåg att de hade stora hunky ögonbrynen också, ochde skulle bli arg och äter snögubbe.
		-- Jack Handey, The New Mexican, 1988.

%
Jag ringde mina föräldrar häromkvällen, men jag glömde bort tidsskillnaden.De är fortfarande lever på femtiotalet.
		-- Strange de Jim

%
Jag gjorde några tunga forskning för att vara förberedda för "Mamma, varför ärhimlen blå? "Han frågade mig om svarta hål i rymden.(Det finns ett hål * där *?)Jag urbenade upp att vara redo för "Varför är gräset grönt?"Han ville diskutera naturens näringskedjor.(Ja, låt oss se, det finns ShopRite, Pathmark ...)Jag talade om Choo-Choo tåg.Han talade förbränningsmotorer.(Förbränningsmotorn sa, "Jag tror att jag kan, jag tror att jag kan.")Jag var nöjd med videospel vurm, tänker vi kunde konkurrerasom jämlikar.Han beskrev komplexiteten i mikrochips som behövs för att skapagrafiken.Sedan puberteten slog. Ah, tonåren.Han sa, "Mamma, jag bara inte förstår kvinnor."(Gotcha!)
		-- Betty LiBrizzi, "The Care and Feeding of a Gifted Child"

%
Jag hatar barn. De är så mänskliga.
		-- H. H. Munro

%
Jag vet vad "vårdnad" [av barnen] betyder. "Ge igen." Det är alltförvar organ. Få även med din gamla dam.
		-- Lenny Bruce

%
Jag älskar barn. Speciellt när de gråter - ty då någon tar bort dem.
		-- Nancy Mitford

%
Jag öppnade lådan i min lilla skrivbord och en enda bokstav föll ut, enbrev från min mor, skriven med blyerts, en av hennes sista, med oavslutadeord och en implicit känsla av hennes avgång. Det är så nyfiken: en kanmotstå tårar och "beter sig" mycket bra i de svåraste timmar av sorg. Mendå någon gör dig en trevlig skylt bakom ett fönster ... eller en meddelandenatt en blomma som var i knopp igår plötsligt har blommat ... ellerett brev glider från en låda ... och allt kollapsar.
		-- Letters From Colette

%
Jag säger ya, jag var en ful unge. Jag var så ful att min pappa höll barnensbild som följde med plånboken han köpte.
		-- Rodney Dangerfield

%
Jag berättade för mina barn, "Someday, du har barn i ditt eget." En av dem sade,"Så kommer du."
		-- Rodney Dangerfield

%
Jag brukade tro att jag var ett barn; Nu tror jag att jag är en vuxen - inte på grundJag inte längre göra barnsliga saker, men eftersom de jag kallar vuxna är intemognare än jag.
		-- Rodney Dangerfield

%
Jag föddes eftersom det var en vana i dessa dagar, människor inte vetnågot annat ... Jag var inte ett barn Prodigy, eftersom ett underbarn ärett barn som vet så mycket när det är ett barn som det gör när det växer upp.
		-- Will Rogers

%
Om ett barn retar dig, lugna honom genom att borsta håret. Om detta intefungerar, använd den andra sidan av borsten på den andra änden av barnet.
		-- Will Rogers

%
Om föräldrarna bara skulle inse hur de bar sina barn.
		-- G. B. Shaw

%
Om graviditet var en bok de skulle skära de två sista kapitlen.
		-- Nora Ephron, "Heartburn"

%
Om mycket gamla kommer ihåg, kommer de mycket unga lyssna.
		-- Chief Dan George

%
Om du har aldrig varit hatad av ditt barn, har du aldrig varit en förälder.
		-- Bette Davis

%
Om din mamma visste vad du gör, skulle hon förmodligen hänga huvudet och gråta.
		-- Bette Davis

%
Sinnessjukdom är ärftlig. Du får den från dina barn.
		-- Bette Davis

%
Det är bättre att förbli barnlös än att skaffa en föräldralös.
		-- Bette Davis

%
Det är inte konstigt att folk är så hemskt när de börjar livet som barn.
		-- Kingsley Amis

%
Det är så snart som jag gjort för jag undrar vad jag börjades för.
		-- Epitaph, Cheltenham Churchyard

%
Det måste ha varit någon ogift dåre som sa "Ett barn kan ställa frågoratt en vis man kan inte svara ", eftersom det i varje anständig hus, en brat sombörjar ställa frågor omgående packad i säng.
		-- Arthur Binstead

%
Det kostar nu mer för att roa ett barn än en gång gjorde att utbilda sin far.
		-- Arthur Binstead

%
Det är aldrig för sent att få en lycklig barndom.
		-- Arthur Binstead

%
Barn ljusna alltid upp ett hus; främst genom att lämna lamporna på.
		-- Arthur Binstead

%
Barnen har * _____ aldrig * tagit vägledning från sina föräldrar. Om du kunderesa tillbaka i tiden och observera den ursprungliga primat familjen iursprungliga trädet, skulle du se primater föräldrar skriker på primatertonåring för att sitta runt och tjura hela dagen i stället för jakt efterlarver och bär som pappa primat. Då skulle du se primatertonåring stampa upp till sin gren och slam bladen.
		-- Dave Barry, "Kids Today: They Don't Know Dum Diddly Do"

%
Lies! Alla lögner! Du alla ligger mot mina pojkar!
		-- Ma Barker

%
Livet börjar inte vid tidpunkten för befruktningen eller födelseögonblicket.Det börjar när barnen lämnar hemmet och hunden dör.
		-- Ma Barker

%
Livet är en sexuellt överförbar sjukdom med 100% dödlighet.
		-- Ma Barker

%
Livet är som en blöja - kort och laddad.
		-- Ma Barker

%
Litteratur är mestadels om att ha sex och inte mycket om att ha barn.Livet är tvärtom.
		-- David Lodge, "The British Museum is Falling Down"

%
Löptid är bara en kort paus i tonåren.
		-- Jules Feiffer

%
Må ni har många vackra och lydiga döttrar.
		-- Jules Feiffer

%
Må ni har många vackra och lydiga söner.
		-- Jules Feiffer

%
Minnen av min familj möten fortfarande är en källa till styrka för mig. jagminns vi hade alla komma in i bilen - jag glömma vilken typ det var - ochköra och köra.Jag är inte säker där vi skulle gå, men jag tror att det fanns några bin där. Delukten av något var stark i luften som vi spelade oavsett sport vispelas. Jag minns en större, äldre kille som vi kallade "pappa". Vi skulle ätavissa saker eller inte och sedan jag tror att vi åkte hem.Jag antar att vissa saker aldrig lämna dig.
		-- Jack Handey, The New Mexican, 1988.

%
Mikrovågor frizz din arvinge.
		-- Jack Handey, The New Mexican, 1988.

%
Min pojke är en genomsnittlig barn. Jag kom hem häromdagen och såg honom tejpa maskartill trottoaren, sitter han där och ser fåglarna få bråck. Väl,bara förra julen jag gav honom en B-B pistol och han gav mig en tröja meden fullträff på baksidan.Jag berättade för mina barn, "Someday, du har barn i ditt eget." En av demsa, "så kommer du."
		-- Rodney Dangerfield

%
Min familj historia börjar med mig, men din slutar med dig.
		-- Iphicrates

%
Min mamma älskade barn - hon skulle ha gett något om jag hade varit en.
		-- Groucho Marx

%
Min mamma sa en gång till mig, "Elwood" (hon alltid kallade mig Elwood)"Elwood, i den här världen du måste vara ack så smart eller ack så trevlig."För år försökte jag smart. Jag rekommenderar trevlig.
		-- Elwood P. Dowde, "Harvey"

%
Min mamma vill barnbarn, så jag sa, "Mamma, go for it!"
		-- Sue Murphy

%
Min mor var ett provrör, min far var en kniv.
		-- Friday

%
Mina föräldrar gick till Niagara Falls och allt jag fick var denna crummy liv.
		-- Friday

%
Min ritual skiljer sig något. Vad jag gör, första [på morgonen], är jaghop i duschkabin. Då jag hop strax tillbaka, eftersom när jag hoppadei jag landade barfota ovanpå See Threepio, lite plast robotkaraktär från "Star Wars" som min son, Robert, gillar att dra benen avav medan han duschar. Sen hoppa tillbaka in i båset, eftersom vår hund,Allvar, som har varit ensam i källaren hela natten bygga upp kraftfullahund känslor, har kommit begränsningsramen och darrande i badrummet och villatt hälsa på mig med 60 eller 70 tusen lekfulla nyp, varav vilken som helst - björni åtanke att jag är naken och utan mina linser i huvudsak blinda- Kan leda till den typ av skada som man måste lära sig en helt nydel om du vill sjunga "Messias", om du får min drivgarn. Då jag hopstrax tillbaka, eftersom Robert, med det kuslig sjätte sinne vissa barnhar - du kan inte lära ut det; de antingen har det eller de inte - har valtexakt det ögonblicket att spola en av toaletterna. Kanske flera av dem.
		-- Dave Barry

%
Natur gör pojkar och flickor vacker att titta på, så att de kan varatolereras tills de får någon mening.
		-- William Phelps

%
har aldrig barn, bara barnbarn.
		-- Gore Vidal

%
låna aldrig bilen till någon som du har fött barn.
		-- Erma Bombeck

%
Höj aldrig handen för att dina barn - det lämnar midsectionoskyddad.
		-- Robert Orben

%
Lita aldrig på en barn längre än du kan kasta det.
		-- Robert Orben

%
Inga hus är childproofed om de små darlings är i tvångströjor.
		-- Robert Orben

%
Oavsett hur gammal en mor är, klockor hon sina medelålders barn förtecken på förbättring.
		-- Florida Scott-Maxwell

%
Ingen lider smärtan av förlossningen eller ångest av att älska ett barn förför presidenter att göra krig, för regeringar att livnära sig på innehållet ideras folk, för försäkringsbolag att lura unga och råna gamla.
		-- Lewis Lapham

%
En far är mer än hundra schoolmasters.
		-- George Herbert

%
En av nackdelarna med att ha barn är att de så småningom blir gamlatillräckligt för att ge dig presenterar de gör i skolan.
		-- Robert Byrne

%
Endast vuxna har svårt med barnsäkra lock.
		-- Robert Byrne

%
Ur munnarna av babes gör ofta kommer spannmål.
		-- Robert Byrne

%
Föräldrar talar ofta om den yngre generationen som om de inte harmycket av något att göra med det.
		-- Robert Byrne

%
Snälla, Mamma! Jag vill hellre göra det själv!
		-- Robert Byrne

%
Reinhart var aldrig hans mors favorit - och han var enda barnet.
		-- Thomas Berger

%
Kom ihåg att som en tonåring du befinner dig i den sista etappen i ditt liv närdu kommer att vara glad att höra att telefonen är för dig.
		-- Fran Lebowitz, "Social Studies"

%
Snö och tonåren är de enda problem som försvinner om du ignorerardem tillräckligt länge.
		-- Fran Lebowitz, "Social Studies"

%
Någonstans på denna jord, var tionde sekund, det är en kvinna som födertill ett barn. Hon måste hittas och stoppas.
		-- Sam Levenson

%
Lär barnen att vara artig och tillmötesgående i hemmet, och när de växer upp,de inte kommer att kunna i kant en bil på en motorväg.
		-- Sam Levenson

%
Provrörs barn bör inte kasta sten.
		-- Sam Levenson

%
Att alla män ska vara bröder är drömmen för människor som inte har några bröder.
		-- Charles Chincholles, "Pensees de tout le monde"

%
Den genomsnittliga inkomsten för den moderna tonåring är cirka 02:00
		-- Charles Chincholles, "Pensees de tout le monde"

%
Rättssalen var gravid (pun intended) med ängslig tystnad somdomare ansåg högtid sin dom i paternitykostym framför honom.Plötsligt nådde han i veck hans kläder, drog ut en cigarr ochhögtid gav den till den tilltalade."Grattis!" deklamerade juristen. "Du har precis blivit enfar!"
		-- Charles Chincholles, "Pensees de tout le monde"

%
Uppsägning av de unga är en nödvändig del av hygien äldremänniskor, och kraftigt hjälper i blodcirkulationen.
		-- Logan Pearsall Smith

%
Det faktum att pojkar tillåts existera alls är ett bevis på en anmärkningsvärdChristian tålamod bland män.
		-- Ambrose Bierce

%
Den första halvan av våra liv är förstört av våra föräldrar och den andra halvanav våra barn.
		-- Clarence Darrow

%
Den fulla effekten av föräldraskap inte slå dig tills du multipliceraAntalet dina barn med trettiotvå tänder.
		-- Clarence Darrow

%
Framtiden är en myt skapad av försäkringsbolag försäljare och high school rådgivare.
		-- Clarence Darrow

%
De goda dör unga - eftersom de ser det är ingen idé att leva om du haratt vara bra.
		-- John Barrymore

%
Tanken är att dö ung så sent som möjligt.
		-- Ashley Montague

%
Den moderna barn kommer att svara dig tillbaka innan du har sagt något.
		-- Laurence J. Peter

%
"Det enda riktiga sättet att se yngre är inte att födas så snart."		   Om och om igen"
		-- Charles Schulz, "Things I've Had to Learn Over and

%
Problemet med genpoolen är att det finns ingen badvakt.
		-- Charles Schulz, "Things I've Had to Learn Over and

%
Det verkliga skälet stora familjer gynna samhället är att åtminstonenågra av barnen i världen bör inte höjas med nybörjare.
		-- Charles Schulz, "Things I've Had to Learn Over and

%
Åren av topp mental aktivitet är utan tvekan i åldrarna fyraoch arton. Vid fyra vi vet alla frågor, vid arton alla svaren.
		-- Charles Schulz, "Things I've Had to Learn Over and

%
"Det var en pojke som heter Eustace Clarence Scrubb, och han nästan förtjänade det."
		-- C. S. Lewis, "The Chronicles of Narnia"

%
Det finns ingen mening med att odlas upp om du inte kan vara barnslig ibland.
		-- Dr. Who

%
Det är inget fel med tonåringar detta resonemang med dem kommer inte att förvärra.
		-- Dr. Who

%
Småbarn är stormtrupper av Lord of Entropy.
		-- Dr. Who

%
Problem är som spädbarn; de bara växa med omvårdnad.
		-- Dr. Who

%
Två moder droppar tillbringade månader att lära sin son hur man ska vara en del avhav. Efter månader av träning, fadern droppen kommenterade till modern droppe,"Vi har lärt vår pojke allt vi vet, han passar att vara tidvattnet."
		-- Dr. Who

%
Vi är alla födda charmig, frisk och spontan och måste vara civiliseradeinnan vi är lämpliga att delta i samhället.Korrekt Behaviour "
		-- Judith Martin, "Miss Manners' Guide to Excruciatingly

%
Vi är människor våra föräldrar varnade oss.
		-- Judith Martin, "Miss Manners' Guide to Excruciatingly

%
Vad som verkligen formar och villkor och gör oss är någon bara ett fåtal avoss någonsin har modet att möta, och det är det barn som du en gång var,långt innan den formella utbildningen någonsin fick sina klor i dig - attotålig, alla krävande barn som vill ha kärlek och kraft och kan inte fånog av endera och som går på rasar och gråtande i din ande tilläntligen ögonen är stängda och alla dårar säga, "Inte han serfredlig? "Det är de uppdämt, sugen barn som gör alla krigoch alla fasor och all konst och all den skönhet och upptäckt iliv, eftersom de försöker uppnå vad som låg utanför deras greppinnan de var fem år gammal.
		-- Robertson Davies, "The Rebel Angels"

%
Vad görs för att barn, kommer de att göra för samhället.
		-- Robertson Davies, "The Rebel Angels"

%
När barndomen dör, är dess lik kallas vuxna.
		-- Brian Aldiss

%
När jag var 16, jag trodde att det inte fanns något hopp för min far. Vid tiden var jag20, han hade gjort stora förbättringar.
		-- Brian Aldiss

%
När du föddes, var en stor chans det tar för dig.
		-- Brian Aldiss

%
Varför de kallar det barnvakt när allt du göra är att köra efter dem?
		-- Brian Aldiss

%
Varför inte ha en gammaldags jul för din familj detta år? Precisbild scenen i vardagsrummet på juldagens morgon som dina barnöppna sina gammaldags presenter.Din 11-åriga son: "Vad sjutton är det här?"Du: "En snurra du snurrar runt, och sedan så småningom fallerner. Vad roligt! Ha, ha! "Son: "Är detta ett skämt Jason Thompson föräldrar fick honom en dator med?två hårddiskar och 128 kilobyte RAM-minne, och jag får dettacretin TOP? "Din 8-åriga dotter: "Du tror att det är illa Titta på den här?".Du: "Det är figgy pudding What a treat!"Dotter: "Det ser ut som get barf."
		-- Dave Barry, "Simple, Homespun Gifts"

%
Du kan lära sig många saker från barn. Hur mycket tålamod du har,till exempel.
		-- Franklin P. Jones

%
"Du kan inte förvänta sig en mamma att vara med ett litet barn hela tiden," MargaretMead anmärkte en gång, med sin vanliga sunt förnuft, men i 1978 hon chockadefeminister genom att snäppa att kvinnor egentligen inte har barn att sätta dem idagvård tolv timmar om dagen, antingen.
		-- Caroline Bird, "The Two Paycheck Marriage"

%
Du kan inte krama ett barn med kärnvapen.
		-- Caroline Bird, "The Two Paycheck Marriage"

%
Ditt ansvar som förälder är inte så stor som man kan föreställa sig. Dubehöver inte förse världen med nästa erövrare sjukdom eller större rörelsebild stjärna. Om ditt barn växer helt enkelt upp att vara någon som inte använderordet "samlar" som ett substantiv, kan du anser dig en okvalificeradframgång.
		-- Fran Lebowitz, "Social Studies"

%
Ungdom är en sådan underbar sak. Vad ett brott att slösa bort den på barn.
		-- George Bernard Shaw

%
Ungdom är förvaltaren av eftervärlden.
		-- George Bernard Shaw

%
Ungdom är när du skylla alla dina bekymmer på era föräldrar; löptidnär du lär dig att allt är fel av den yngre generationen.
		-- George Bernard Shaw

%
Ungdom. Det är ett under att någon någonsin outgrows det.
		-- George Bernard Shaw

%
