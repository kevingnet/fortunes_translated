En tysk, en stolpe och en tjeckisk vänster läger för en vandring genom skogen.Efter att ha rapporterades saknad en dag eller två senare, rangers hittade två björnar,en en hane, en kvinnlig, ser misstänkt overstuffed. de dödadehonan, obducerades henne, och att det finns tillräckligt fann tyska och polacken.	"Vad tror du?" sade den första ranger."Den tjeckiska är i den manliga", svarade den andra.
		-- Guindon

%
Aberdeen var så liten att när familjen med bilen gickpå semester, bensinstationen och drive-in teater var tvungna att stänga.
		-- Guindon

%
Enligt Rand McNally platser rankade almanacka, det bästa stället att bo iAmerika är staden Pittsburgh. Staden New York kom i tjugofemte.Här i New York vi verkligen inte bryr sig för mycket. Eftersom vi vet att vi kundeslå upp sin stad som helst.
		-- David Letterman

%
"Alla ormar som vill stanna kvar i Irland kommer att glädja höja deras högra hand."
		-- Saint Patrick

%
Dessutom är skottarna sägs ha uppfunnit golf. Då hade deatt uppfinna skotsk whisky för att ta bort smärtan och frustration.
		-- Saint Patrick

%
alta, v: För att ändra; göra eller bli annorlunda; ändra.Ansa, V: a talat eller skriftligt svar, som på en fråga.baa, N: a plats människor träffas för att ha ett par drinkar.Baaston, n: huvudstad Massachusetts.baaba, n: En vars verksamhet är att klippa eller trimma hår eller skägg.beea, n: En alkoholhaltig dryck bryggs från malt och humle, oftahittas i baas.caaa, n: En bil.Centa, n: En punkt kring vilken något kretsar; axel. (Ellernågon som arbetar med Knicks.)chouda, n: En tjock skaldjurssoppa, ofta i en mjölk bas.dada, n: Information, esp. information som organiseras för analys ellerberäkning.
		-- Massachewsetts Unabridged Dictionary

%
Amerika upptäcktes av Amerigo Vespucci och namngavs efter honom, tillsmänniskor fick trötta på att leva i en plats som heter "Vespuccia" och byttenamn till "Amerika".
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Amerika, hur kan jag skriva en helig litania i fåniga humör?
		-- Allen Ginsberg

%
Amerikan vid födelse; Texan vid nåden av guden.
		-- Allen Ginsberg

%
Amerikaner är människor som insisterar på att leva i nuet, spänd.
		-- Allen Ginsberg

%
Amerikanernas största rädsla är att Amerika kommer att visa sig ha varit enfenomen, inte en civilisation.
		-- Shirley Hazzard, "Transit of Venus"

%
En amerikansk är en man med två armar och fyra hjul.
		-- A Chinese child

%
En engelsman har aldrig själv, med undantag för ett ädelt syfte.
		-- A. P. Herbert

%
Allt någon kan säga om Amerika är sant.
		-- Emmett Grogan

%
Armenier och azerier i Stepanakert, huvudstad i Nagorno-Karabachautonoma regionen, upplopp över välbehövlig stavningsreformen i Sovjetunionen.
		-- P. J. O'Rourke

%
Baseball är en skicklig spel. Det är USA: s spel - det, och höga skatter.
		-- The Best of Will Rogers

%
Bond återspeglas att goda amerikaner var fina människor och att de flesta av demtycktes komma från Texas.
		-- Ian Fleming, "Casino Royale"

%
Boston State House är navet i solsystemet. Du kan inte bända ut detav en Boston man om du hade däcket i hela skapelsen rätas ut för enkofot.
		-- Oliver Wendell Holmes

%
Carol huvud värkte när hon släpade bakom unsmiling Calibreeslängs block av bås. Hon chirruped på Kennicott, "Låt oss vara vild!Låt oss rida på Merry-go-round och ta en guldring! "Kennicott ansåg det, och mumlade att Calibree, "Tänk dig folksvill stoppa och prova en åktur på Merry-go-round? "Calibree ansåg det, och mumlade till sin hustru, "Tror du att du villatt stoppa och prova en åktur på Merry-go-round? "Fru Calibree log i en urtvättad sätt, och suckade, "Åh nej,Jag tror inte jag bryr mig för mycket, men du folks gå vidare och prova det. "Calibree uppges Kennicott, "Nej, jag tror inte att vi bryr oss till enhel del, men du folks gå vidare och prova det. "Kennicott sammanfattade hela målet mot vildhet: "Låt oss försökadet en annan gång, Carrie. "Hon gav upp.
		-- Sinclair Lewis, "Main Street"

%
Klimat och kirurgiR C Gilchrist, som sköts av J Sharp tolv dagar sedan, och somfick en derringer boll i höger bröst, och som det var tänkt påtiden kan inte leva flera timmar, var på gatan i går ochdagen före - gå flera block samtidigt. Till dem som utformar att varafull av kulor eller skurna i bitar med Bowie-knivar, vi hjärtligtrekommenderar vår Sacramento klimat och Sacramento kirurgi.
		-- Sacramento Daily Union, September 11, 1861

%
David Letterman s "Saker som vi kan vara stolta över som amerikaner":* Största antalet medborgare som faktiskt har bordade ett UFO* Många tidningar funktionen "RÖRA"* timma motell* De allra flesta Elvis filmer görs här* Inte bara ge upp direkt under andra världskrigetsom vissa länder vi kan nämna* Goatees & Van Dykes tros endast bäras av weenies* Våra skötsam golfproffs* Fabulous babes kust till kust
		-- Sacramento Daily Union, September 11, 1861

%
Decemba, n: Den 12: e månaden på året.erra, n: Ett misstag.faa, n: till, från eller på betydande avstånd.Linder, n: En kvinnlig namn.Memba, n: För att hämta till sinnet; tänka på igen.New Hampsha, n: en stat i nordöstra USA.New Yaak, n: en annan stat i nordöstra USA.Novemba, n: Den 11: e månaden på året.Octoba, n: Den 10: e månaden på året.ägg, n: Location ovanför eller över en viss position. Vad isäsongen är när Knicks sluta spela.
		-- Massachewsetts Unabridged Dictionary

%
Detroit är Cleveland utan glitter.
		-- Massachewsetts Unabridged Dictionary

%
Gör Miami en tjänst. När du lämnar, ta någon med dig.
		-- Massachewsetts Unabridged Dictionary

%
Vet du Montana?
		-- Massachewsetts Unabridged Dictionary

%
Vet du skillnaden mellan en yankee och en damyankee?En yankee kommer söderut till * _____ besök *.
		-- Massachewsetts Unabridged Dictionary

%
Eli och Bessie gick att sova.Mitt i natten, Bessie puffade Eli."Var så vänlig och stänga fönstret. Det är kallt ute!"Halvsovande, mumlade Eli,"Nu ... så om jag ska stänga fönstret, kommer det att vara varmt ute?"
		-- Massachewsetts Unabridged Dictionary

%
Fem personer - en engelsman, ryska, amerikanska, fransman och Irishmanvar och ombedd att skriva en bok om elefanter. Viss tid senare dealla hade avslutat sina respektive böcker. Engelsmannen bok hade rätt"The Elephant - Hur att samla in dem", den ryska "The Elephant -. Vol I",den amerikanska "The Elephant - Hur man tjäna pengar på dem", fransmannens"The Elephant - dess parning vanor" och irländaren "The Elephant ochIrländsk politisk historia ".
		-- Massachewsetts Unabridged Dictionary

%
Av någon anledning passerar en glasyr över människors ansikten när du säger"Kanada". Vi kanske borde invadera South Dakota eller något.
		-- Sandra Gotlieb, wife of the Canadian ambassador to the U.S.

%
Fortune presenterar:Användbara fraser på esperanto # 1.^ Cu VI parolas vinkel? Pratar du engelska?Mi ne komprenas. jag förstår inte.Vi estas la sola esperantisto kiun mi Du är den enda Esperanto högtalarerenkontas. Jag har träffat.La ^ Ceko estas enpo ^ stigita. Kontrollen är i posten.Oni ne povas, ^ gin netrovi. Du kan inte missa det.Mi nur rigardadas. Jag tittar bara.Nu, ^ sajnis bona ideo. Tja, det verkade som en bra idé.
		-- Sandra Gotlieb, wife of the Canadian ambassador to the U.S.

%
Fortune presenterar:Användbara fraser på esperanto # 2.^ Cu tiu loko estas okupita? Är den här platsen upptagen?^ Cu vi ofte Venas ^ ci-tien? Kommer du hit ofta?^ Cu mi povas havi via telelonnumeron? Kan jag få ditt telefonnummer?Mi estas komputilisto. Jag jobbar med datorer.Mi legas multe da scienca fikcio. Jag läser en hel del science fiction.^ Cu necesas ke vi eliras? Har du verkligen att gå?
		-- Sandra Gotlieb, wife of the Canadian ambassador to the U.S.

%
Fortune presenterar:Användbara fraser på esperanto # 5.Mi ^ cevalovipus vin se mi havus Jag skulle hästpiska dig om jag hade en häst.^ Cevalon.Vere VI ^ sercas. Skojar du.Nu, parDOOOOOnu min! Tja exCUUUUUSE mig!Kiu invitis vin? Som bjuder in dig?Kion vi diris pri mia Patrino? Vad sa du om min mamma?Bu ^ så ^ stopu min per kulero. Gag mig med en sked.
		-- Sandra Gotlieb, wife of the Canadian ambassador to the U.S.

%
Gay shlafen: Yiddish för "somna".Nu inte "gay shlafen" har en mjukare, mer lugnande ljud än denhårda, staccato "somnar"? Lyssna på skillnaden:"Gå att sova, du lilla stackare!" ... "Gay shlafen, älskling."Självklart, är inte det?Klart det bästa du kan göra för dig barn är att börjatalar jiddisch just nu och aldrig tala ett ord i engelska somlänge du lever. Detta kommer naturligtvis att innebära undervisning Jiddisch till alladina vänner, affärsbekanta, folk i snabbköpet, ochså vidare, men det är bara poängen. Det måste börja med engageradeindivider och sedan växa ....Vissa mindre justeringar måste göras, naturligtvis: detecken skrivna i vad ser ut Yiddish bokstäver kommer inte att vara roligt närallt är skrivet på jiddisch. Och vi måste börja köra påden vänstra sidan av vägen så att vi inte kommer att läsa gatuskyltarbakåt. Men är det ett alltför högt pris att betala för världsfreden?Jag tror inte, min vän, jag tror inte det.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
"Gee, Toto, jag tror inte att vi är i Kansas längre."
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
"Gud ger bördor, också axlar"Jimmy Carter citerade denna judiska talesätt i sitt koncessions tal vidslutet av 1980 valet. Åtminstone sade han att det var en judisk talesätt; jagkan inte hitta det någonstans. Jag är säker på att han talar sanning men; varförskulle han ljuga om något sådant?
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
God natt, Austin, Texas, var du än är!
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Hating Yankees är som amerikan som pizza paj, ogifta mödrar ochfusk på din inkomstskatt.
		-- Mike Royko

%
Har du sett den senaste japanska kamera? Tydligen är det så fort det kanfotografera en amerikansk med munnen stängd!
		-- Mike Royko

%
Hör om den kaliforniska terrorist som försökte spränga en buss?Brände läpparna på avgasröret.
		-- Mike Royko

%
Hör om den unga kinesiska kvinnan som just vunnit på lotto?En lyckosam kaka ...
		-- Mike Royko

%
Här är det faktum att veckan, kanske till och med det faktum att i månaden.Enligt förmodligen tillförlitliga källor, är Coca-Cola människor uppleversvår marknadsföring ångest i Kina.Orden "Coca-Cola" översätta till kinesiska som antingen (beroendepå böjnings) "vax-göds mare" eller "bita vaxet grodyngel".Bita vaxet grodyngel.Det finns ett slags grov rättvisa, är det inte?Problemet med detta faktum, så vacker som den är, är att det är svårtatt få en hel kolumn av det. Jag skulle vilja lära världen att bita ett vaxgrodyngel. Coke - det är den verkliga vax-göds sto. Inte illa, men bredsatiric perspektiv när inte öppna upp.
		-- John Carrol, The San Francisco Chronicle

%
"Hans stora mål var att fly från civilisationen, och så snart han hadepengar, gick han till södra Kalifornien. "
		-- John Carrol, The San Francisco Chronicle

%
Historiker har nu definitivt fastställts att Juan Cabrillo, upptäckKalifornien, inte var ute efter Kansas, vilket skapar ett prejudikat somfortsätter än i dag.
		-- Wayne Shannon

%
Houdini flyr från New Jersey!Film på elva.
		-- Wayne Shannon

%
Hur många präster behövs för en Boston Mass?
		-- Wayne Shannon

%
Jag är bara en fin, ren skuren mongoliska pojke.
		-- Yul Brynner, 1956

%
Jag är, i själva verket, en särskilt hotfulla och exklusiv person, avpre-Adamite ancestral härkomst. Du kommer att förstå detta när jag berättaatt jag kan spåra min anor tillbaka till en protoplasmal ursprunglig atommetallkorn. Därför är min familj stolthet något otänkbart. jagkan inte hjälpa det. Jag föddes hånfull.
		-- Pooh-Bah, "The Mikado"

%
Jag visste inte att han var död; Jag trodde att han var brittisk.
		-- Pooh-Bah, "The Mikado"

%
Jag har definierat hundra procent amerikan som nittionio procent en idiot.
		-- George Bernard Shaw

%
Jag sköt en pil in i luften, och det fastnade.På en klar dag,U.C.L.A.Det finns så mycket föroreningar i luften nu att om det inte vore för vårlungor det skulle finnas någon plats att sätta allt.
		-- Robert Orben

%
Jag går igenom min "Jag vill gå tillbaka till New York" fas idag. händervarje halvår eller så. Så tänkte jag, kanske oklokt att jag skulle deladen med dig.> I New York i vintern är det miljoner minusgrader och  vinden färdas på en miljon miles i timmen ner 5th avenue.> Och i LA är det 72.> I New York i sommaren är det en miljon grader och luftfuktigheten  är en miljon procent.> Och i LA är det 72.> I New York finns det en miljon intressanta människor.> Och i LA finns 72.
		-- Robert Orben

%
"Jag är i Pittsburgh. Varför är jag här?"
		-- Harold Urey, Nobel Laureate

%
Om alla kinesiska samtidigt hoppade i Stilla havet utanför en 10 fotplattform uppfördes 10 fot utanför deras kust, skulle det orsaka en flodvågsom skulle förstöra allt i det här landet väster om Nebraska.
		-- Harold Urey, Nobel Laureate

%
Illinois är inte precis det land som Gud glömde - det är mer somland Han försöker ignorera.
		-- Harold Urey, Nobel Laureate

%
År 1880 den franska fångade Detroit men gav det tillbaka ... de kunde intefå delar.
		-- Harold Urey, Nobel Laureate

%
I Amerika, det är inte hur mycket en artikelkostnader, det är hur mycket du sparar.
		-- Harold Urey, Nobel Laureate

%
I alla världens menyn, måste Kanada anses vara vichyssoise nationer -det är kallt, halv-franska, och svårt att röra.
		-- Stuart Keate

%
I Kalifornien de inte kasta sina sopor bort - de gör det iTV-program.
		-- Woody Allen, "Annie Hall"

%
I Minnesota frågar de varför alla fotbollsplaner i Iowa har konstgräs.Det är så cheerleaders inte betar under spelets gång.
		-- Woody Allen, "Annie Hall"

%
Indiana är ett tillstånd tillägnad basket. Basket, sojabönor, svin ochbasketboll. Berkeley, onödigt att säga, är inte alls lika atletisk. Berkeleyär tillägnad kaffe, ångest, gropar och kaffe.
		-- Carolyn Jones

%
Inglish Spocken Hier: några sargade översättningarLogga på en hyttdörr av en sovjetisk Svarta havet kryssningsfartyget:Helpsavering apparata i emergings si många visselpipor!Koppla strängarna apparata om bosums och träffabakom, flyr sedan till likgiltig lifesaveringshippenobedicing de instruerar i kärlet.På dörren i ett hotell i Belgrad:Låt oss veta om någon unficiency samt läcker ut på		tjänsten. Vårt yttersta kommer att förbättra den.
		-- Colin Bowles

%
Inglish Spocken Hier: några sargade översättningarLogga på en katedral i Spanien:Det är förbjudet att ange en kvinna, även en utlänning omklädd som en man.Ovanför enterance till en Kairo bar:Ensamkommande damer inte medgav inte med makeeller liknande.På Bukarest hiss:Hissen är fastställs för de kommande dagarna.Under den tiden beklagar vi att du kommer att vara outhärdligt.
		-- Colin Bowles

%
Inglish Spocken Hier: några sargade översättningarOlika tecken i Polen:Högersväng mot omedelbar utanför.Gå lugnande i snön, eftersom det lurar skid demoner.Fem o'clock tea på alla timmar.I en för män toalett i Sidney:Skaka överflödigt vatten från händer, tryck knappen för att starta,gnugga händerna snabbt under luftuttaget och torka händernapå framsidan av skjortan.
		-- Colin Bowles, San Francisco Chronicle

%
Iowans frågar varför Minnesotans inte dricka mer Kool-Aid. Det är för attde kan inte räkna ut hur man får två liter vatten i en av demsmå papperskuvert.
		-- Colin Bowles, San Francisco Chronicle

%
Är inte det trevligt att människor som föredrar Los Angeles till San Francisco bor där?
		-- Herb Caen

%
Det är svårt att hävda att Gud hatade Oklahoma. Om han inte gjorde det, varför är det sånära Texas?
		-- Herb Caen

%
Det är inte Camelot, men det är inte Cleveland, heller.
		-- Kevin White, Mayor of Boston

%
Det räcker inte med att vara ungersk; du måste ha talang också.
		-- Alexander Korda

%
Det är märkligt och lite oroande, att reflektera över det faktum attEngelska är det enda större språk som "I" aktiveras; i mångaandra språk "Du" aktiveras och "jag" är gemener.
		-- Sydney J. Harris

%
Det är egentligen ganska enkelt val: liv, död, eller Los Angeles.
		-- Sydney J. Harris

%
Att lära sig franska är trivialt: ordet för hästen är cheval, och allt annatföljer på samma sätt.
		-- Alan J. Perlis

%
Som så många amerikaner, hon försöker bygga ett liv som gjordekänsla av saker som hon hittade i presentbutiker.
		-- Kurt Vonnegut, Jr.

%
Likaså nationella aptitretare, saltlösning cured sill med rå lök,vinner några vänner, undantaget tyskarna.
		-- Darwin Porter "Scandinavia On $50 A Day"

%
Att bo i LA är som att inte ha ett datum på lördag kväll.
		-- Candice Bergen

%
Bor i New York ger människor verkliga incitament att vilja saker somingen annan vill.
		-- Andy Warhol

%
Minnesota -hem för blont hår och blå öron.mygga leverantör till den fria världen.kommer att bli kär i en lom.där besökarna blir blå med avund.en dag det är varmt, resten av året det är kallt.land med många kulturer - mestadels i halsen.där eliten träffas slask.handske it or leave it.många är kallt, men få är frysta.land av skidan och hem för galna.mark 10.000 Peter.
		-- Andy Warhol

%
Moishe Margolies, som vägde hela 105 pounds och stod en ännu fem foti hans strumpor, tog sin första flygplan resa. Han tog plats bredvid enklumpig bruiser av en man som råkade vara tungviktvärlden. Little Moishe var orolig nog innan han ens kom in i planet,men nu bruset av motorer och den stora höjden absolut livrädd honom.Så rädd blev han att hans mage vänds och han kastade upp alltöver muskel jätte lokaliseringen bredvid honom. Lyckligtvis, åtminstone för Moishe,Mannen var god sömn. Men nu den lille mannen hade ett annat problem. how ivärlden skulle han någonsin förklara situationen till bastant brute när hanvaknat? Den plötsliga röst värdinna på planets intercom slutligenvaknade bruiser och Moishe, hans hjärta i hans mun, ökade till tillfälle."Känsla bättre nu?" frågade han solicitously.
		-- Andy Warhol

%
Monterey ... är avgjort mest trivsamma och mest civiliserade utseende platsi Kalifornien ... [det] är också en utmärkt plats för kuk-fighting, spelav olika slag, Fandangos, och olika typer av nöjen och knavery.
		-- Richard Henry Dama, "Two Years Before the Mast", 1840

%
De flesta Texans tror Hanukkah är något slags anka samtal.
		-- Richard Lewis

%
Mina godda välsigna, aldrig ser jag Sucha människor.
		-- Signor Piozzi, quoted by Cecilia Thrale

%
New York är verklig. Resten görs med speglar.
		-- Signor Piozzi, quoted by Cecilia Thrale

%
New York leder nu världens stora städer i antalet människor runtsom du inte bör göra en plötslig rörelse.
		-- David Letterman

%
Oavsett vilka andra nationer kan säga om USA,invandring är fortfarande den ärligaste formen av smicker.
		-- David Letterman

%
"Och Herren Gud planterade en trädgård öster om Whittier på en plats som heterYorba Linda, och ur marken han gjorde att odla apelsinträd somvar bra för mat och frukterna därav han märkt SUNKIST ... "
		-- "The Begatting of a President"

%
På natten innan hennes familj flyttade från Kansas till Kalifornien, den lillaflicka knäböjde vid sin säng att säga hennes böner. "Gud välsigne mamma och pappa ochKeith och Kim ", sade hon. När hon började att stiga upp, hon snabbt till," Åh,och Gud, är detta adjö. Vi flyttar till Hollywood. "
		-- "The Begatting of a President"

%
På det hela taget, skulle jag hellre vara i Philadelphia.
		-- W. C. Fields' epitaph

%
En av reglerna för Busmanship, New York stil, aldrig ge upp dinsäte till en annan passagerare. Detta kan verka känslolöst, men det är det bästasätt, verkligen. Om en passagerare skulle ge en plats till någon som svimmadei gången, säg, de andra på bussen skulle bli förvirrad ochföreställa sig att de var i Topeka Kansas.
		-- W. C. Fields' epitaph

%
paak, n: en arena eller inclosed spelplan. Att sätta eller lämna (enett fordon) för en tid i en viss plats.patato, n: stärkelse, ätbara knöl av en allmänt odlad växt.Septemba, n: Den 9: e månaden på året.Sua, n: Har ingen tvekan; viss.sista, n: En kvinnlig med samma mor och far som högtalaren.Tamato, n: en köttig, slätskaliga rödaktig frukt äts i salladereller som en grönsak.Troopa, n: En stat polis.Wista, n: En stad i centrala Masschewsetts.yaad, n: ett område av marken intill en byggnad.
		-- Massachewsetts Unabridged Dictionary

%
Kanske, trots allt, Amerika aldrig har upptäckts. Jag själv skullesäger att det bara hade upptäckts.
		-- Oscar Wilde

%
Philadelphia är inte tråkig - det bara verkar så eftersom det är bredvidspännande Camden, New Jersey.
		-- Oscar Wilde

%
Providence, New Jersey, är en av de få städer där Velveeta ostvisas på gourmet hyllan.
		-- Oscar Wilde

%
San Francisco är inte vad det brukade vara, och det var aldrig.
		-- Herb Caen

%
Seattle är så våt att människor skydda sin egendom med watch-ankor.
		-- Herb Caen

%
Verkar att en opinionsundersökare tog en global opinionsundersökning.Hennes fråga var, "Ursäkta mig, Vad är din åsikt om köttbrist"I Texas, svaret var "Vad är en brist?"I Polen, svaret var "Vad är kött?"I Sovjetunionen, var svaret "Vad är en åsikt?"I New York, var svaret "Vad är ursäkta mig?"
		-- Herb Caen

%
Vissa 1500 miles väster om Big Apple finner vi Minneapple, enoas av lugn i oroliga tider. Det är en bra stad, en civiliserad stad.En stad där de fortfarande vet hur man får dina skjortor tillbaka genom torsdag. LåtaBig Apple har bedrifter av "Broadway Joe" Namath. Vi har känttröga men stadig Killebrew. Lyssna på Cole Porter över en dry martinikan mycket väl passa dem otur aldrig har hört Whoopee John PolkaBand och aldrig har delat en kanna 3,2 Grain Belt öl. Förlusten ärderas. Och Big Apple har ännu inte baka bagel som kan matcha jordnötsmör på lefse. Här är en stad där den viktiga urban problemet är holländska almsjukdom och antalet ett brott är övertidsparkering. Vi skryter mer teaterper capita än Big Apple. Vi går att se, inte ses. Vi går ävennär vi måste skyffla tio inches av snö från uppfarten för att komma dit. Verkligenvintrarna är hård. Men sedan kommer förundras av Minneapple sommaren.Folk flockas till stadens sjöar att leka och glädjas vid åsynen av såmycket glad mänskligheten fri från bindningar av den traditionella ned fyllda parkas.Här finns till Minneapple. Och dess folk. Vår känsla för stil är balanseradgenom en hälsosam respekt för vind chill faktorer.Och vi alltid, alltid äta våra grönsaker.Detta är den Minneapple.
		-- Herb Caen

%
Någon gjorde en studie av de tre mest ofta hört fraser i New YorkStad. Den ena är "Hej, taxi." Två är "Vad tåg tar jag för att komma tillBloomingdales? "Och tre är," Var inte orolig. Det är bara ett köttsår. "
		-- David Letterman

%
"Någonstans", sa fader Vittorini, "gav Blake inte tala omMaskinerier av glädje? Det vill säga, inte Gud främja miljöer, dåskrämma dessa naturer genom provocera förekomsten av kött, leksaks män ochkvinnor, såsom är vi alla? Och så glatt sänt ut, på vårt bästa, medbra nåd och fina intelligens, på lugna Noons, i verkligt klimat, är vi inte GudsMaskinerier av glädje? ""Om Blake sade att", sa fader Brian "han bodde aldrig i Dublin."
		-- R. Bradbury, "The Machineries of Joy"

%
Den Allsmäktige i sin oändliga vishet såg inte lämpligt att skapa fransmäni bilden av engelsmännen.
		-- Winston Churchill, 1942

%
Den amerikanska nationen i den sjätte avdelningen är en fin folk; de älskareagle - på baksidan av en dollar.
		-- Finlay Peter Dunne

%
Den anglosaxiska samvete hindrar inte anglosaxiska frånSinning, bara hindrar det honom från att njuta av sin synd.
		-- Salvador De Madariaga

%
I bästa fall: Få lön från Amerika, bygga ett hus i England,leva med en japansk hustru, och äta kinesisk mat.Ganska bra fall: Få lön från England, bygga ett hus i Amerika,leva med en kinesisk fru, och äta japansk mat.Det värsta fallet: Få lön från Kina, bygga ett hus i Japan,leva med en brittisk fru och äta amerikansk mat.
		-- Bungei Shunju, a popular Japanese magazine

%
Det bästa som kommer ut ur Iowa är I-80.
		-- Bungei Shunju, a popular Japanese magazine

%
De stora städerna i Amerika blir länder i tredje världen.
		-- Nora Ephron

%
Britterna kommer! Britterna kommer!
		-- Nora Ephron

%
Klimatet i Bombay är sådant att invånarna måste bo någon annanstans.
		-- Nora Ephron

%
Förbannelse irländska är inte att de inte vet orden till en sång -det är att de känner dem * ___ alla *.
		-- Susan Dooley

%
Tjeckerna meddelade efter Sputnik att de också skulle starta en satellit.Naturligtvis skulle det bana Sputnik, inte jorden!
		-- Susan Dooley

%
Skillnaden mellan USA och England är att engelska tror 100miles är en lång sträcka och amerikanerna tror 100 år är en lång tid.
		-- Susan Dooley

%
Ägget grädde är psykologiskt motsatsen till omskärelse - det* Pleasurably * bekräftar din judiskhet.
		-- Mel Brooks

%
Den engelska godsägare galopperande efter en räv - det outsägligafullt driva kvickhuvud.
		-- Oscar Wilde, "A Woman of No Importance"

%
Den engelska har ingen respekt för deras språk, och kommer inte att lärasina barn att tala det.
		-- G. B. Shaw

%
Den engelska instinktivt beundrar någon människa som inte har någon talang och är blygsamom det.
		-- James Agate, British film and drama critic

%
[Den franska Rivieran är] en solig plats för skumma människor.
		-- Somerset Maugham

%
Den geografiska centrum Boston är i Roxbury. På grund norr omcentrum finner vi den södra änden. Detta är inte att förväxla med SouthBoston som ligger direkt öster om South End. Norr om SouthEnd är East Boston och sydväst om East Boston är norra ände.
		-- Somerset Maugham

%
De goys har visat följande sats ...föreläsning.
		-- Physicist John von Neumann, at the start of a classroom

%
Mars landade hans tefat på Manhattan, och omedelbart efterväxande blev kontaktad av en panhandler. "Mister", sade mannen, "kan jaghar en fjärdedel? "Mars frågade: "Vad är en fjärdedel?"Den panhandler tänkte en minut, lyste, sedan sa, "Du ärhöger! Kan jag har en dollar? "
		-- Physicist John von Neumann, at the start of a classroom

%
Den mygga är den statliga fågeln av New Jersey.
		-- Andy Warhol

%
Det vanligaste tilltalsnamn i världen är Mohammad; den vanligasteefternamn i världen är Chang. Kan ni föreställa er det enorma antaletmänniskor i världen som heter Mohammad Chang?
		-- Derek Wills

%
Den enda kulturella fördelen LA har över NY är att du kan göra en rättaktivera ett rött ljus.
		-- Woody Allen

%
San Diego Freeway. Officiell parkeringen av 1984 OS!
		-- Woody Allen

%
Problemet är, det finns ett oändligt utbud av vita Män, men det haralltid varit ett begränsat antal människohandel.
		-- Little Big Man

%
Världens mest ivrig baseboll fan (en Aggie) hade kommit tillstadion för det första spelet i World Series bara att inse att han hade lämnathans biljett hemma. Inte vill missa något av den första omgången, gick hantill biljettluckan och fick i en lång rad för en annan sits. Efter en timmesvänta han var bara ett par fötter från montern när en röst ropade, "Hey,Dave! "The Aggie såg upp, klev ut ur linje och försökte hitta ägarenav rösten - utan framgång. Sedan insåg han att han hade förlorat sin plats ilinje och fick vänta över igen. När fläkten slutligen köpte sin biljett,han var törstig, så han gick för att köpa en drink. Linjen vid koncession montervar lång, också, men eftersom spelet inte hade började han bestämde sig för att vänta. Precis somHan kom till fönstret, en så kallad röst, "Hej, Dave!" Återigen Aggie försöktatt hitta rösten - men ingen lycka. Han var mycket upprörd när han kom tillbaka i linjeför hans drink. Slutligen fan gick till sin plats, ivriga för spelet att börja.När han väntade på planen, hörde han röstsamtal, "Hey Dave!" en gång till.Rasande, stod han upp och skrek på toppen av sina lungor, "Mitt namn är inte Dave!"
		-- Little Big Man

%
Sedan fanns det Formosan bartendern som heter Taiwan-On.
		-- Little Big Man

%
Det * __ är * intelligent liv på jorden, men jag lämnar för Texas på måndagen.
		-- Little Big Man

%
Det finns människor som tycker att det är konstigt att äta fyra eller fem kinesiska måltiderpå rad; i Kina, jag påminna dem ofta, det finns en miljard eller såmänniskor som tycker inget konstigt om det.
		-- Calvin Trillin

%
Det är inget fel med södra Kalifornien som en ökning avhavsytan skulle inte bota.
		-- Ross MacDonald

%
Det måste finnas minst 500.000.000 råttor i USA; självklart,Jag har aldrig hört historien förut.
		-- Ross MacDonald

%
Det var en gång denna swami som bodde över en delicatessan. verkar endag bestämde han att stanna i bottenvåningen för lite frisk lever. Jo, ägareav deli var lite av en billig-skridsko, och bestämde sig för att plocka upp lite extraändra på sin kundens bekostnad. Turning tyst till counterman, hanviskade: "tynga på swami lever!"
		-- Ross MacDonald

%
Det var en New Yorker som hade en livslång ambition att vara en Texan.Lyckligtvis hade han en Texan vän och gick till honom för att få råd. "Mikrofon,du vet att jag har alltid velat vara en Texan. Du är en * ____ verklig * Texan, vadborde jag?""Jo", svarade Mike, "Det första du måste göra är att sesom en Texan. Det innebär att du måste klä rätt. Den andra sakendu har att göra är att tala i en sydlig drawl. ""Tack, Mike, jag ska ge det ett försök," svarade New Yorker.Några veckor gått och New Yorker släntrar in i en butik kläddi en tio-liters hatt, cowboykängor, Levi jeans och en bandana. "Hallå där,pardner, jag vill ha lite nötkött, inte alltför sällsynta, och vissa av dem färska kex, "Han berättar counterman.Killen bakom disken tar en lång titt på honom och sedan säger,"Du måste vara från New York."New Yorker rodnar, och säger: "Ja, ja, jag är. Hur gjordedu vet?""Eftersom detta är en järnaffär."
		-- Ross MacDonald

%
Det är bara något jag inte tycker om Virginia; staten.
		-- Ross MacDonald

%
Det är något annorlunda med oss ​​- skiljer sig från människor i Europa,Afrika, Asien ... en djup och varaktig tro på påskharen.
		-- G. Gordon Liddy

%
Tre Midwesterners, en Kansan, en Missourian och en Iowan,allt som förekommer på ett frågesportprogram, ombads att fylla i den här meningen:"Gamla MacDonald hade en...""Gamla MacDonald hade en förgasare," svarade Kansan."Tyvärr, det är fel," spelet programledare sa."Gamla MacDonald hade en broms justering nedåt påbensinstation ", sade Missourian."Fel"."Gamla MacDonald hade en gård", sade Iowan.	"KORREKT!" ropar quizmaster. "Nu för $ 100.000, stava" gård ".""Easy", sade Iowan. "E-I-E-I-O."
		-- G. Gordon Liddy

%
Tippa över hela världen på sin sida och allt löst kommer att landa i Los Angeles.
		-- Frank Lloyd Wright

%
Till en kalifornisk, måste en person visa sig kriminellt sinnessjuka innan hantillåts att köra taxi i New York. För New York cabbies, ärlighet ochstannar vid rött ljus är båda tillval.
		-- From "East vs. West: The War Between the Coasts

%
Till en kalifornisk, alla New York-bor är kallt; även i värme de sällan gåröver femtioåtta grader. Om du kollapsar på en gata i New York, planatt tillbringa några dagar där.
		-- From "East vs. West: The War Between the Coasts

%
Till en New Yorker, alla kalifornier är blond, även de svarta. Det finns,i själva verket hela stadsdelar som är planlagd endast för blonda personer. Deenda sättet att skilja mellan Kalifornien och Sverige är att denSvenskarna talar bättre engelska. "
		-- From "East vs. West: The War Between the Coasts

%
Till en New Yorker, de enda Kalifornien hus på marknaden för mindre än enmiljon dollar är de i brand. Dessa går i allmänhet för sexhundratusen.
		-- From "East vs. West: The War Between the Coasts

%
För att vara lycklig man måste vara a) väl utfodras, unhounded av simpla bekymmer, till mods iZion, b) full av en behaglig känsla av överlägsenhet till massorna av ensandra män, och c) fint och oupphörligt roade enligt en smak.Det är min uppfattning att om denna definition godtas, finns det inget landi världen där en man bildade som jag - en man med min säregnasvagheter, fåfänglighet, aptit och aversioner - kan vara så glad som han kanvara i USA. Going vidare, jag fastställa doktrinen att det ären ren fysisk omöjlighet för en sådan människa att leva i USAoch inte vara glad.
		-- H. L. Mencken, "On Being An American"

%
Att veta Edina är att förkasta det.
		-- Dudley Riggs, "The Year the Grinch Stole the Election"

%
Toto, jag tror inte att vi är i Kansas anymore.
		-- Judy Garland, "Wizard of Oz"

%
Turister - ha lite kul med New Yorks hårdkokta cabbies. När dukomma till din destination, säg till din förare, "Betala? Jag var liftade."
		-- David Letterman

%
Trafiksignaler i New York är bara grova riktlinjer.
		-- David Letterman

%
Reser genom New England, en bilist stannade för gas i en liten by."Vad är det här ställe som heter?" frågade han stationen skötare."Allt beror," de infödda drawled. "Menar du med dem som haratt leva i denna pappa-skulden, malätna, damm täckta, en-hoss dumpa, ellerav dem som är bara att njuta av dess pittoreska och pittoreska rustika charmför ett kort pass? "
		-- David Letterman

%
Besök vackra Vergas, Minnesota.
		-- David Letterman

%
Besök vackra Wisconsin Dells.
		-- David Letterman

%
Besök [1] den vackra Smoky Mountains![1] besök, v .:Kom för en vecka, spendera för mycket pengar och betala massor av dolda skatter,sedan lämna. Vi ska vara glada att se dina pengar igen nästa år.Du kan spara tid genom att helt enkelt skicka pengar, om du är för upptagen.
		-- David Letterman

%
Vi bryr oss inte hur de gör det i New York.
		-- David Letterman

%
Välkommen till Lake Wobegon, där alla män är starka, kvinnorna är vackra,och barnen är över genomsnittet.
		-- Garrison Keillor

%
Vilken typ av smutsiga affärer är du på nu? Jag menar, man ditgår du? Vart går du, Amerika, i din glänsande bil på natten?
		-- Jack Kerouac

%
Oavsett inte lyckas i två månader och en halv i Kalifornien kommeraldrig lyckas.
		-- Rev. Henry Durant, founder of the University of California

%
När en man är trött på London är han trött på livet.
		-- Samuel Johnson

%
När kommer sommaren kommit till Minnesota, frågar du? Tja, förra året, jagtror att det var en tisdag.
		-- Samuel Johnson

%
När jag först kom i detta land jag hade bara femton cent i fickanoch en vilja att kompromissa.
		-- Weber cartoon caption

%
När jag såg en skylt på motorvägen som sagt, "Los Angeles 445 miles", sa jagför mig själv, "jag måste komma ur denna bana."
		-- Franklyn Ajaye

%
När du vant sig vid att aldrig vara ensam, kan du anser digAmericanized.
		-- Franklyn Ajaye

%
Skulle den sista personen att lämna Michigan vänd ut ljuset?
		-- Franklyn Ajaye

%
Yawd [substantiv, Bostonese]: campus Ha Id.
		-- Webster's Unafraid Dictionary

%
Ja, jag har nu fått denna fina lilla lägenhet i New York, en av demL-formade sådana. Tyvärr är det en gemena l.
		-- Rita Rudner

%
Du har alltid möjlighet att pitching baseballs på tomma sprayburkari en cul-de-sac i en förort till Cleveland.
		-- Rita Rudner

%
Du behöver inte flytta till Edina, du uppnå Edina.
		-- Guindon

%
Du vet att du är i en liten stad vid ...Du behöver inte använda blinkers eftersom alla vet vart du ska.Du är född den 13 juni och din familj får gåvor från lokalahandlarna för att du är det första barnet av året.Alla vet vars kredit är bra, och vars fru är inte.Du talar till varje hund du passerar genom namn ... och han viftar på svansen.Du slår fel nummer, och prata i 15 minuter i alla fall.Du skriver en check på fel bank och det täcker dig ändå.
		-- Guindon

%
