1 tjurar, 3 kor.
		-- Leo Costales, in "Outside July 2005"

%
3000000 $.
		-- Leo Costales, in "Outside July 2005"

%
40 är inte gammal. Om du är ett träd.
		-- Leo Costales, in "Outside July 2005"

%
En galande ligger högst upp sig själv på en telefontråd. Han skulle göra enlångväga caw.
		-- Leo Costales, in "Outside July 2005"

%
En furore Normanorum libera nos, O Domine![Från raseri norsemen befria oss, o Herre!]
		-- Medieval prayer

%
En logg kan flyta i en flod, men det gör inte det en krokodil.
		-- Medieval prayer

%
En pickup med tre killar i den drar in i lumber varvet. En av de mänkommer ut och går in på kontoret."Jag behöver ungefär fyra-by-två-talet", säger han."Du måste betyda två och fyra s" svarar expediten.Mannen repor huvudet. "Vänta en minut", säger han, "jag ska gåkolla upp."Tillbaka efter en animerad konversation med andra passagerare ilastbil, försäkrar han expediten att, ja, i själva verket, två och fyra skulle varagodtagbar."OK", säger expediten, skriva ner det, "hur länge du vill ha dem?"Killen får tom blick igen. "Öh ... Jag antar att jag bättre gåkontrollera ", säger han.Han går tillbaka till lastbilen, och det finns en annan animeradkonversation. Killen kommer tillbaka till kontoret. "En lång tid", säger han,"Vi bygger ett hus".
		-- Medieval prayer

%
En förutsägelse är värd tjugo förklaringar.
		-- K. Brecher

%
En vördnads ville ringa en annan vördnads. Han berättade operatören,"Detta är en parson att parson samtalet."
		-- K. Brecher

%
En gummiskrapa med något annat namn skulle inte låta som roligt.
		-- K. Brecher

%
Ett vakuum är en fan så mycket bättre än några av de saker som naturenersätter det med.
		-- Tennessee Williams

%
En ung flicka, Carmen Cohen, kallades av hennes efternamn av sin far,och hennes första namn av sin mor. När hon var tio, inte visste om honvar Carmen eller Cohen.
		-- Tennessee Williams

%
Enligt min bästa minne, jag minns inte.
		-- Vincent "Jimmy Blue Eyes" Alo

%
Vuxna dör ung.
		-- Vincent "Jimmy Blue Eyes" Alo

%
African Violet: En sådan värd är sällsyntÄppelblom: preferensKandidat knapp: CelibatLagerblad: Jag förändras, men i dödenCamelia: Reflekterad DezereKrysantemum, röd: Jag älskarKrysantemum, vit: SanningenKrysantemum, andra: förolämpat kärlekKlöver: Var minCrocus: Abuse intePåsklilja: InnocenceFörgätmigej inte: Sann kärlekFuchsia: SnabbGardenia: Secret, outsägligt kärlekKaprifol: band av kärlekIvy: Vänskap, trohet, äktenskapJasmine: Amiablity, transporter av glädje, sensualitetLöv (döda): MelancholyLila: Ungdomlig oskuldLilly: Renhet, sötmaLilly av dalen: Return of lyckaMagnolia: Värdighet, uthållighet* En upp-och-ned blossom reverserar betydelsen.
		-- Vincent "Jimmy Blue Eyes" Alo

%
Ålder är en tyrann som förbjuder vid straff i livet, alla njutningar av ungdomar.
		-- Vincent "Jimmy Blue Eyes" Alo

%
Håller med dem nu, det kommer att spara så mycket tid.
		-- Vincent "Jimmy Blue Eyes" Alo

%
Ah, tsarens basar bisarra beaux-arts!
		-- Vincent "Jimmy Blue Eyes" Alo

%
Ahhhhhh ... lukten av Cuprinol och mahogny. Det retar mig att ...handlingar av passion ... handlingar ... oduglighet.
		-- Vincent "Jimmy Blue Eyes" Alo

%
Alla telefonsamtal är oanständigt.
		-- Karen Elizabeth Gordon

%
Alla riktigt bra idéer som jag någonsin haft kom till mig medan jag mjölka en ko.
		-- Grant Wood

%
Jag påfluget? Jag hoppas det. Min påfluget blir raves.
		-- Grant Wood

%
Fantastiskt men sant ...Om allt lax fångad i Kanada under ett år lades ände till ändeöver Saharaöknen, skulle lukten vara helt fruktansvärt.
		-- Grant Wood

%
Fantastiskt men sant ...Det finns så mycket sand i norra Afrika som om det spreds ut detskulle helt täcka Saharaöknen.
		-- Grant Wood

%
Amnesia brukade vara min favorit ord, men då jag glömde det.
		-- Grant Wood

%
En atom-blaster är ett bra vapen, men det kan peka åt båda hållen.
		-- Isaac Asimov

%
... Och dessutom ... Jag gillar inte dina byxor.
		-- Isaac Asimov

%
Och jag ensam är återvände till vifta på svansen.
		-- Isaac Asimov

%
Någon sten i start vandrar alltid mot tryckgradienten tillexakt den punkt där de flesta tryck.
		-- Milt Barber

%
Varje gång saker och ting verkar gå bättre, har du missat något.
		-- Milt Barber

%
Är vi inte män?
		-- Milt Barber

%
Som Zeus sade till Narcissus, "Titta på dig själv."
		-- Milt Barber

%
Avec!
		-- Milt Barber

%
BAD vansinne MAN !!!
		-- Milt Barber

%
Barfota magnetisera vassa metallföremål så att de pekar uppåt frångolv - särskilt i mörker.
		-- Milt Barber

%
Batterier ingår ej.
		-- Milt Barber

%
VAR UPPMÄRKSAM!!!! (Världen behöver fler lerts ...)
		-- Milt Barber

%
VARA BORTA! (Det har varit en ny befolkningsexplosion av lerts.)
		-- Milt Barber

%
Innan jag visste den bästa delen av mitt liv hade kommit, hade det gått.
		-- Milt Barber

%
Bli frustrerade är obehaglig, men de verkliga katastrofer i livet börjarnär du får vad du vill.
		-- Milt Barber

%
Tro allt du hör om i världen; ingenting är alltför omöjligt dåligt.
		-- Honor'e de Balzac

%
Största säkerhets gap - en öppen mun.
		-- Honor'e de Balzac

%
Bizarreness är kärnan i det exotiska.
		-- Honor'e de Balzac

%
Skyll Saint Andreas - det är hans fel.
		-- Honor'e de Balzac

%
Välsignade är de som går runt i cirklar, ty de skall kallas Wheels.
		-- Honor'e de Balzac

%
Blå färg idag.[Roligt Jack Slingwine, Guy Harris och Hal Pierson. Ed.]
		-- Honor'e de Balzac

%
Pojke! Eukalyptus!
		-- Honor'e de Balzac

%
Pojke, som krita säker gjorde ont!
		-- Honor'e de Balzac

%
Bushydo - vägen för buske. Bonsai!
		-- Honor'e de Balzac

%
"Men Huey, du lovade!""Säg att jag ljög."
		-- Honor'e de Balzac

%
Men i likhet med bibeln säger ... Det finns större affärer framöver!
		-- Honor'e de Balzac

%
Av uthållighet snigeln nådde Ark.
		-- Charles Spurgeon

%
CF & C stal det, rättvist och torg.
		-- Tim Hahn

%
Kapitel VIIIPå grund av konvergensen av krafter bortom hans fattningsförmåga, SalvatoreQuanucci plötsligt sprutade ut ur universum som en vattenmelonfrö, och aldrig hört från igen.
		-- Tim Hahn

%
Färglösa gröna idéer sova ursinnigt.
		-- Tim Hahn

%
Confucius något att säga för mycket.
		-- Recent Chinese Proverb

%
Grattis är i ordning för Tom Reid.Han säger att han fick just reda på att han är vinnaren av 2021 psykiska avYear.
		-- Recent Chinese Proverb

%
Kultur är vana att bli nöjd med det bästa och att veta varför.
		-- Recent Chinese Proverb

%
Custer begått Siouxicide.
		-- Recent Chinese Proverb

%
"Oavsett saknade massan i universum är, jag hoppas att det inte kackerlackor!"
		-- Mom

%
Död åt alla fanatiker!
		-- Mom

%
Avgår i bitar, det vill säga, split.
		-- Mom

%
Beröva en spegel av sitt silver och även tsaren kommer inte se hans ansikte.
		-- Mom

%
Sa jag två? Jag ljög.
		-- Mom

%
Har det någonsin inträffa för er att fett chans och smal chans betyder samma sak?Eller att vi kör på ways och parkera på uppfarter?
		-- Mom

%
Hörde du om modellen som satt på en trasig flaska och skär en fin siffra?
		-- Mom

%
Visste du ...Att ingen någonsin läser dessa saker?
		-- Mom

%
"Die? Jag skulle säga inte, käre vän. Ingen Barrymore skulle tillåta en sådankonventionell sak att hända honom. "
		-- John Barrymore's dying words

%
Värdighet är som en flagga. Den flaxar i en storm.
		-- Roy Mengot

%
Dime är pengar.
		-- Roy Mengot

%
Inte underskatta kraften i Force.
		-- Roy Mengot

%
Använd inte det främmande ord "ideal". Vi har det bra inföddaordet "lögner".
		-- Henrik Ibsen, "The Wild Duck"

%
Tycker folk vet att du har fräknar överallt?
		-- Henrik Ibsen, "The Wild Duck"

%
Tycker eleverna i Zenbuddism do Om-arbete?
		-- Henrik Ibsen, "The Wild Duck"

%
"Tror du på intuition?""Nej, men jag har en konstig känsla av att jag en dag kommer."
		-- Henrik Ibsen, "The Wild Duck"

%
Har du lysdexia?
		-- Henrik Ibsen, "The Wild Duck"

%
Har du försonande socialt värde?
		-- Henrik Ibsen, "The Wild Duck"

%
Har en enbent anka simma i en cirkel?
		-- Henrik Ibsen, "The Wild Duck"

%
Tvinga inte, få en större hammare.
		-- Anthony

%
Inte gissa - kontrollera dina säkerhetsbestämmelser.
		-- Anthony

%
Inte jag vet att du?
		-- Anthony

%
Låt inte din status blir alltför quo!
		-- Anthony

%
Sluta inte nu, kan vi lika gärna låsa dörren och kasta bort nyckeln.
		-- Anthony

%
Inte tala om tid, tills du har talat med honom.
		-- Anthony

%
Oroa dig inte - det brontosaurus är långsam, dum, och lugn.
		-- Anthony

%
Oroa dig inte om du är en kleptoman; du kan alltid ta något för det.
		-- Anthony

%
Dubbel!
		-- Anthony

%
Dr Jekyll hade något Hyde.
		-- Anthony

%
Dr Livingston?Dr Living I. förmodar?
		-- Anthony

%
Rita på min fina kommando av språket, sa jag ingenting.
		-- Anthony

%
Drömmar är gratis, men det finns en liten avgift för ändringar.
		-- Anthony

%
Släppa att pickle!
		-- Anthony

%
Släpp vas och det kommer att bli en Ming av det förflutna.
		-- The Adventurer

%
Duckies är kul!
		-- The Adventurer

%
Ankor? Vad ankor ??
		-- The Adventurer

%
Dungeons & Dragons är bara en massa Saxon våld.
		-- The Adventurer

%
Under ett slagsmål, en man kastade en skål med Jello på sin hustru. Hon hadehonom arresterad för att bära ett stelnat vapen.I en annan kamp, ​​hustru dekorerad honom med en tung glaskanna.Hon är en kvinna som conks att dvala.
		-- The Adventurer

%
Dyslexi innebär aldrig behöva säga att du är ysror.
		-- The Adventurer

%
Dyslexics har mer FNU.
		-- The Adventurer

%
Dyslexics av ​​världen, UNTIE!
		-- The Adventurer

%
"Jorden är en stor, stor funhouse utan kul."
		-- Jeff Berner

%
Redigering är en omformulering aktivitet.
		-- Jeff Berner

%
Eggheads förena er! Du har inget att förlora, men dina äggulor.
		-- Adlai Stevenson

%
Händelser påverkas inte, utvecklar de.
		-- Sri Aurobindo

%
Någonsin undrar varför brandbilar är röda?Eftersom tidningar läses också.Två och två är fyra.Fyra och fyra är åtta.Åtta och fyra är tolv.Det finns tolv inches i en linjal.Queen Mary var en linjal.Queen Mary var ett skepp.Fartygen seglar havet.Det finns fiskar i havet.Fiskar har fenor.Finländarna slogs ryssarna.Ryssarna är röda.Brandbilar är alltid Rush'n.Därför brandbilar är röda.
		-- Sri Aurobindo

%
Varje absurditet har en mästare som kommer att försvara den.
		-- Sri Aurobindo

%
Varje dag är det samma sak - sort. Jag vill ha något annorlunda.
		-- Sri Aurobindo

%
Varje gång jag tror att jag vet var det är på, de flyttar den.
		-- Sri Aurobindo

%
Varje gång du lyckas stänga dörren på verkligheten, det kommer in genomfönster.
		-- Sri Aurobindo

%
Varje ord är som en onödig fläck på tystnad och intet.
		-- Beckett

%
Allt bågar till framgång, även grammatik.
		-- Beckett

%
Allt kan göras under "diverse".
		-- Beckett

%
Allt kan vara olika i detta om bara en sak hadevarit annorlunda i det förflutna.
		-- Beckett

%
Allt ska byggas top-down, utom den första gången.
		-- Beckett

%
Allt ska byggas top-down, men den här gången.
		-- Beckett

%
Allt tar längre tid, kostar mer och är mindre användbara.
		-- Erwin Tomash

%
Allt du vet är fel!
		-- Erwin Tomash

%
Fakta upphör inte att existera eftersom de ignoreras.
		-- Aldous Huxley

%
Fakta, bortsett från deras relationer, är som etiketter på tomma flaskor.
		-- Sven Italla

%
"Fantasier är gratis.""NEJ !! NEJ !! Det är tankepolisen !!!!"
		-- Sven Italla

%
Långt mattare än en orm tand det är att tillbringa en lugn ungdom.
		-- Sven Italla

%
Fetter Loves Madelyn.
		-- Sven Italla

%
Att ta reda på vad som händer i C.I.A. är som utför akupunkturpå en klippa.
		-- New York Times, Jan. 20, 1981

%
Fem cyklar gör en Volkswagen, sju gör en lastbil.
		-- Adolfo Guzman

%
Flamma!
		-- Johnny Storm

%
Fly mig bort till den ljusa sidan av månen ...
		-- Johnny Storm

%
För en helig stint, en mal av duken gav upp sina ylle för ludd.
		-- Johnny Storm

%
För dig den undergörande jorden sätter fram söta blommor.
		-- Titus Lucretius Carus

%
Tvinga den !!!Om den går sönder, ja, det fungerade inte i alla fall ...Nej, inte tvinga den, få en större hammare.
		-- Titus Lucretius Carus

%
Tvinga dig själv att slappna av!
		-- Titus Lucretius Carus

%
Skogsbränder orsakar Smokey björnar.
		-- Titus Lucretius Carus

%
Fortune graffito i veckan (eller kanske till och med månad):Skriv inte på väggarna!(Och under)Du vill jag ska skriva?
		-- Titus Lucretius Carus

%
Fortune kontor Dörrskylt av veckan:Oförbätterlig VITSMAKARE - inte incorrige.
		-- Titus Lucretius Carus

%
"Fann det" musen svarade ganska vresigt: "naturligtvis du vetvad det betyder.""Jag vet vad det betyder väl nog, när jag hittar en sak", sadeDuck: "det är i allmänhet en groda eller en mask Frågan är, vad gjorde.ärkebiskop hitta? "
		-- Titus Lucretius Carus

%
Från en viss punkt och framåt finns det inte längre någon återvändo.Det är den punkt som måste uppnås.
		-- F. Kafka

%
Rasande aktivitet är ingen ersättning för att förstå.
		-- H. H. Williams

%
Allmänna begrepp är i allmänhet fel.
		-- Lady M. W. Montagu

%
Ge mig en rörmokare vän storleken på Pittsburgh kupolen, och en platsatt stå, och jag kommer att dränera världen.
		-- Lady M. W. Montagu

%
GE UPP!!!!
		-- Lady M. W. Montagu

%
Med tanke på mina druthers, skulle jag druther inte.
		-- Lady M. W. Montagu

%
Gloffing är ett tillstånd av mig.
		-- Lady M. W. Montagu

%
Gå "sätt! Du stör mig!
		-- Lady M. W. Montagu

%
Gå bort, jag är okej.
		-- H. G. Wells' last words.

%
Gå klättra en gravitations väl!
		-- H. G. Wells' last words.

%
Mål ... Planer ... de är fantasier, de är en del av en drömvärld ...
		-- Wally Shawn

%
Gud är död.Nietzsche är död.Nietzsche är Gud.
		-- Dead

%
Gud är inte död, han bara inte kunde hitta en parkeringsplats.
		-- Dead

%
Gud är inte död. Han bara inte vill engagera sig.
		-- Dead

%
Gud skapade världen på sex dagar, och greps på sjunde.
		-- Dead

%
Gud var nöjd med sitt eget arbete, och det är dödlig.
		-- Samuel Butler

%
Gud, jag ber om tålamod - och jag vill ha det just nu!
		-- Samuel Butler

%
Goda nyheter är bara livets sätt att hålla dig ur balans.
		-- Samuel Butler

%
Half Moon i kväll. (Åtminstone är det bättre än ingen månen alls.)
		-- Samuel Butler

%
Lycka gör upp i höjd vad det saknar i längd.
		-- Samuel Butler

%
Glad fest gris!
		-- Samuel Butler

%
Hårda verkligheten har ett sätt att kramper din stil.
		-- Daniel Dennett

%
Har på dig!
		-- Daniel Dennett

%
Ha modet att ta dina egna tankar på allvar, för de kommer att forma dig.
		-- Albert Einstein

%
"Har du bott här hela ditt liv?""Åh, dubbelt så länge."
		-- Albert Einstein

%
Har du låst din arkivskåp?
		-- Albert Einstein

%
Har ni märkt att allt du behöver för att växa frisk, är kraftig gräs enspricka i trottoaren?
		-- Albert Einstein

%
"Han kastade sig på sin häst och red madly i alla riktningar."
		-- Albert Einstein

%
Den som tillbringar en storm under ett träd, tar livet med en nypa TNT.
		-- Albert Einstein

%
Hedonist att hyra ... inget jobb för lätt!
		-- Albert Einstein

%
Hjälp en svala landa på Capistrano.
		-- Albert Einstein

%
Hjälp stämpla ut och avskaffa redundans och upprepning.
		-- Albert Einstein

%
HJÄLP! Man fångade i en människokropp!
		-- Albert Einstein

%
HJÄLP! Skrivmaskinen är bruten!
		-- E. E. CUMMINGS

%
Här det finnas tygers.
		-- E. E. CUMMINGS

%
"Hans ögon var kall. Så kallt som den bittra vintern snö som föllutanför. Ja, kall och därför svår att tugga ... "
		-- E. E. CUMMINGS

%
Tuta, om du hatar bildekaler som säger "Tuta om ..."
		-- E. E. CUMMINGS

%
Tuta, om du älskar lugn och ro.
		-- E. E. CUMMINGS

%
Hushållsarbete kan döda dig om det görs rätt.
		-- Erma Bombeck

%
Hur kan du vara på två ställen på en gång när du inte någonstans alls?
		-- Erma Bombeck

%
Hur kommer det bara dina vänner steg på din nya vita sneakers?
		-- Erma Bombeck

%
Hur kommer det sig att vi aldrig prata längre?
		-- Erma Bombeck

%
Hur kommer fel nummer är aldrig upptagen?
		-- Erma Bombeck

%
Hur snällt av dig att vara villiga att leva någons liv för dem.
		-- Erma Bombeck

%
Hur mycket av sitt inflytande på dig är ett resultat av ditt inflytande på dem?
		-- Erma Bombeck

%
Hur untasteful kan du få?
		-- Erma Bombeck

%
Va?
		-- Erma Bombeck

%
Jag vaknar alltid upp i crack i is.
		-- Joe E. Lewis

%
Jag är mor till allt, och allt ska bära en tröja.
		-- Joe E. Lewis

%
Jag kan läsa dina tankar, och du bör skämmas.
		-- Joe E. Lewis

%
Jag kan relatera till det.
		-- Joe E. Lewis

%
Jag kan motstå allt annat än frestelsen.
		-- Joe E. Lewis

%
Jag kunde omöjligen undgå att hålla med dig mindre.
		-- Joe E. Lewis

%
Jag föraktar nöjet att tilltalande människor som jag föraktar.
		-- Joe E. Lewis

%
Jag har inte någon lösning, men jag beundrar verkligen problemet.
		-- Ashleigh Brilliant

%
"Jag har inget emot att gå ingenstans så länge det är en intressant väg."
		-- Ronald Mabbitt

%
Jag förstår dig inte längre.
		-- Ronald Mabbitt

%
Jag vill inte att synas alltför nyfikna, men är du fortfarande lever?
		-- Ronald Mabbitt

%
Jag tycker den tid som vi tillbringar tillsammans.
		-- Ronald Mabbitt

%
Jag existerar, därför är jag betalat.
		-- Ronald Mabbitt

%
Jag är rädd förklaringar förklarande saker förklaras.
		-- Ronald Mabbitt

%
Jag tycker synd om din hjärna ... ensam i den stora stort huvud ...
		-- Ronald Mabbitt

%
"Jag fick reda på varför min bil humming. Det hade glömt orden."
		-- Ronald Mabbitt

%
Jag hatar citat.
		-- Ralph Waldo Emerson

%
Jag hatar troll. Kanske kunde jag Metamorph det till något annat - som englupande, två huvuden, eldsprutande drake.
		-- Willow

%
Jag har en fruktansvärd huvudvärk, jag var att sätta på toaletten vatten och locket föll.
		-- Willow

%
Jag har blivit mig utan mitt samtycke.
		-- Willow

%
Jag har fler träffpunkter som du möjligt kan tänka dig.
		-- Willow

%
Jag har sett den stora Pretender och han är inte vad han verkar.
		-- Willow

%
Jag har inte förlorat mitt sinne; Jag vet exakt var jag lämnade det.
		-- Willow

%
Jag hör ljudet att maskinerna gör och känna mitt hjärta paus, baraför ett ögonblick.
		-- Willow

%
Jag hör vad du säger, men jag bryr mig inte.
		-- Willow

%
Jag vet allt. Jag kan bara inte komma ihåg allt på en gång.
		-- Willow

%
Jag vet att du tror att du trodde att du visste vad du trodde jag sa,men jag är inte säker på att du förstått vad du trodde jag menade.
		-- Willow

%
Jag vet att du är på jakt efter sig själv, jag bara inte har sett dig någonstans.
		-- Willow

%
Jag lever som jag skriver; snabb, med en hel del misstag.
		-- Willow

%
Jag älskar förräderi men hatar en förrädare.
		-- Gaius Julius Caesar

%
Jag gjorde aldrig det sättet förut.
		-- Gaius Julius Caesar

%
"Jag rör bara bas med verkligheten på ett behov när det behövs!"
		-- Royal Floyd Mengot (Klaus)

%
[Jag tänker] för att se, höra, röra, och förstöra allt i min väg,inklusive rödbetor, kålrötter, och mest slumpmässiga grönsaker, men med undantag av jams,som jag absolut livrädd för jams ...Egentligen tror jag att min rädsla för jams började i min tidiga ungdom, då mångaav mina unga kamrater bombarderade mig med detsamma för att sjunga sånger av fjärran länderoch djupa blå hav på ett språk i hög grad liknar den hos den gemensamma suggan.Min psykos var ytterligare imponerade i min själ som jag nått tonåren,när, medan hoppa genom ett fält av jams, lättsamt gungade blommori stratosfären, slet en stor yam-picking maskin genom fälten,förfölja mig till kanten av den stora plantage, där jag flydde genom att dykatill ett stort dike fylls med en blandning av vatten och svingödsel, vilket kanförklara min tendens att skrika, "Här kommer mars! Göm äggen!" varjetid jag har fläsk. Men jag göra en utvikning. Faktum kvarstår att jag kan inte rationelltitu med jams, och grisar är fruktansvärda conversationalists.
		-- Royal Floyd Mengot (Klaus)

%
Jag förutspår att i dag kommer att bli ihåg förrän i morgon!
		-- Royal Floyd Mengot (Klaus)

%
Jag vägrar att ha en kamp om förstånd med en obeväpnad person.
		-- Royal Floyd Mengot (Klaus)

%
Jag såg vad du gjorde och jag vet vem du är.
		-- Royal Floyd Mengot (Klaus)

%
Jag luktar Wumpus.
		-- Royal Floyd Mengot (Klaus)

%
Jag trodde att du tystade vakten!
		-- Royal Floyd Mengot (Klaus)

%
Jag förstår varför du är förvirrad. Du tänker för mycket.
		-- Carole Wallach.

%
Jag brukade vara en agnostiker, men nu är jag inte så säker.
		-- Carole Wallach.

%
Jag brukade få hög på livet, men på sistone har jag byggt upp ett motstånd.
		-- Carole Wallach.

%
Jag brukade tro att jag var obeslutsamma, men nu är jag inte så säker.
		-- Carole Wallach.

%
Jag vill nå dig - där det för närvarande ligger?
		-- Carole Wallach.

%
Jag kommer alltid att älska den falska bild jag hade av dig.
		-- Carole Wallach.

%
Jag kommer att göra dig kortare vid huvudet.
		-- Elizabeth I

%
Jag kommer aldrig att ljuga för dig.
		-- Elizabeth I

%
Jag kommer inte att glömma dig.
		-- Elizabeth I

%
Jag skulle inte vara så paranoid om du inte var allt för att få mig !!
		-- Elizabeth I

%
Jag skulle vara en sämre människa om jag aldrig hade sett en örn fluga.[Jag såg en örn flyga en gång. Lyckligtvis hade jag min eagle flugsmälla praktiskt. Ed.]
		-- John Denver

%
Jag skulle ge min högra arm att vara ambidextrous.
		-- John Denver

%
"Jag dör" han kraxade."Min experiment var en succé," kemisten svarade."Du kan inte riktigt träna en beagle," han dogmatiserat."Det är ingen beagle, det är en blandras" muttrade hon."Elden går ut", han vrålade."Dålig skytte," jägaren groused."Du borde se en psykiater," han påminde mig."Du orm" hon skramlade."Någon är vid dörren," hon instämde."Bolagets kommande", säger hon gissade."Dawn kom för tidigt", säger hon sörjde."Jag tror att jag ska avsluta det hela," Sue suckade."Jag beställde choklad, inte vanilj," Jag skrek."Din broderi är slarvig" hon nålade grymt."Var har du fått detta kött?" han tyglad hest.
		-- Gyles Brandreth, "The Joy of Lex"

%
Jag är glad att jag inte är född före te.
		-- Sidney Smith (1771-1845)

%
Jag kommer att ta upp en fråga och hålla den i örat.
		-- John Foreman

%
Jag skrattar inte med dig, jag skrattar åt dig.
		-- John Foreman

%
Jag är inte erbjuda mig själv som ett exempel; varje liv utvecklas genom sina egna lagar.
		-- John Foreman

%
Jag är inte fördomsfull, jag hatar alla lika.
		-- John Foreman

%
Jag är inte stolt.
		-- John Foreman

%
Jag är inte spänd, bara hemskt, fruktansvärt alert!
		-- John Foreman

%
Jag är beredd för alla nödsituationer men helt oförberedd för det dagliga livet.
		-- John Foreman

%
Jag är så bröt jag kan inte ens uppmärksamma.
		-- John Foreman

%
Jag har flyttats!
		-- John Foreman

%
Jag har varit där.
		-- John Foreman

%
Jag har haft ungefär lika mycket av detta som jag kan stå.
		-- John Foreman

%
Identifiera dina besökare.
		-- John Foreman

%
Lättja är en resa för dårar.
		-- John Foreman

%
"Om en kamel flugor, skrattar ingen om det inte blir mycket långt."
		-- Paul White

%
Om alla män var bröder, skulle du låta en gifta din syster?
		-- Paul White

%
Om allt kommer din väg då är du i fel körfält.
		-- Paul White

%
Om allt verkar gå bra, har du uppenbarligen förbisett något.
		-- Paul White

%
Om Gud är död, som kommer att rädda drottningen?
		-- Paul White

%
Om Gud är en, vad är dåligt?
		-- Charles Manson

%
Om jag kunde släppa död just nu, skulle jag vara den lyckligaste mannen vid liv!
		-- Samuel Goldwyn

%
Om jag inte ser dig i framtiden, jag ser dig i hagen.
		-- Samuel Goldwyn

%
Om jag älskar dig, vilken verksamhet är det din?
		-- Johann van Goethe

%
Om det inte luktar ännu, är det ganska färskt.
		-- Dave Johnson, on dead seagulls

%
Om det häller före sju, har det regnat av elva.
		-- Dave Johnson, on dead seagulls

%
Om det inte var så varmt i dag, skulle det vara svalare.
		-- Dave Johnson, on dead seagulls

%
Om det inte vore för den sista minuten, skulle ingenting någonsin blir gjort.
		-- Dave Johnson, on dead seagulls

%
Om livet ger dig citroner, gör lemonad.
		-- Dave Johnson, on dead seagulls

%
Om livet är bara ett skämt, fortfarande kvarstår frågan: för vars nöjen?
		-- Dave Johnson, on dead seagulls

%
Om livet är inte vad du ville, du har bett om något annat?
		-- Dave Johnson, on dead seagulls

%
Om kaniner fötter är så lyckliga, vad hände med kaninen?
		-- Dave Johnson, on dead seagulls

%
Om ändarna inte helgar medlen, vad gör?
		-- Robert Moses

%
Om det engelska språket gjorde någon mening, skulle kompromissar ha någotatt göra med en brist på blommor.[För att inte nämna, fjäril vore flutterby. Ed.]
		-- Doug Larson

%
Om framtiden är inte vad det brukade vara, betyder det att det förflutnakan komma att ändras i tider framöver?
		-- Doug Larson

%
Om gräset är grönare på andra sidan staketet, överväga vad som kan varafertilizing den.
		-- Doug Larson

%
Om betydelsen av "sant" och "falskt" har bytt, då denna meningskulle inte vara falsk.
		-- Doug Larson

%
Om oddsen är en miljon till ett mot något inträffar, är chansenär 50-50 det kommer.
		-- Doug Larson

%
Om det inte finns någon Gud, som dyker upp nästa Kleenex?
		-- Art Hoppe

%
Om tiden läker alla sår, hur kommer naveln förblir densamma?
		-- Art Hoppe

%
Om vi ​​ser ljuset i slutet av tunneln, är det mot bakgrund av enmötande tåg.
		-- Robert Lowell

%
Om du ska gå på tunn is, kan man lika gärna dansa.
		-- Robert Lowell

%
Om du kan leda den till vatten och tvinga den att dricka, är det inte en häst.
		-- Robert Lowell

%
Om du inte tänka på framtiden, kan du inte ha en.
		-- John Galsworthy

%
Om du har något att göra, inte göra det här.
		-- John Galsworthy

%
Om du visste vad jag ska säga härnäst, skulle du säga det?
		-- John Galsworthy

%
Om du vet svaret på en fråga, fråga inte.
		-- Petersen Nesbit

%
Om du sticka huvudet i sanden, är en sak säker, du kommerfå din bak sparkas.
		-- Petersen Nesbit

%
Om du är rätt 90% av tiden, varför käbbla om de återstående 3%?
		-- Petersen Nesbit

%
Fantasin sätter ett vapen i kriget mot verkligheten.
		-- Jules de Gaultier

%
Tänk vad vi kan föreställa oss!
		-- Arthur Rubinstein

%
Immanuel inte vits, han Kant.
		-- Arthur Rubinstein

%
Immanuel Kant men Kubla Khan.
		-- Arthur Rubinstein

%
I händelse av brand, står i hallen och ropa "Fire!"
		-- The Kidner Report

%
I min slut är min början.
		-- Mary Stuart, Queen of Scots

%
I kriget om förstånd, han är obeväpnad.
		-- Mary Stuart, Queen of Scots

%
I denna värld, kan sanningen vänta; Hon är van vid det.
		-- Mary Stuart, Queen of Scots

%
Inkludera mig.
		-- Mary Stuart, Queen of Scots

%
Obeslutsamhet är den sanna grunden för flexibilitet.
		-- Mary Stuart, Queen of Scots

%
Likgiltighet kommer säkerligen att vara undergång mänskligheten, men vem bryr sig?
		-- Mary Stuart, Queen of Scots

%
Sömnlöshet är inte något att förlora sömn över.
		-- Mary Stuart, Queen of Scots

%
Är döden rättsligt bindande?
		-- Mary Stuart, Queen of Scots

%
Är inte flygresor underbart? Frukost i London, middag i New York,bagage i Brasilien.
		-- Mary Stuart, Queen of Scots

%
Det har länge varit känt att fåglar emellanåt kommer att bygga bon imanar av hästar. Den enda kända lösningen på detta problem är att ströbagerijäst i manen, för, som vi alla vet, är jäst jäst och boär boet, och aldrig manen ska tweet.
		-- Mary Stuart, Queen of Scots

%
Det är en lärdom som alla historien lär vise män, att sätta tilltro till idéer,och inte under omständigheter.
		-- Emerson

%
Det är bättre att aldrig ha fötts. Men vem av oss har sådan tur?One in a million, kanske.
		-- Emerson

%
Det är bättre att vara hjulbent än ingen ben.
		-- Emerson

%
Det är bättre att kyssa en avokado än att få i ett slagsmål med en jordsvin.
		-- Emerson

%
Det är lättare att motstå i början än vid slutet.
		-- Leonardo da Vinci

%
Det är lättare att köra nedför en backe än upp en.
		-- Leonardo da Vinci

%
Det är verksamheten i framtiden att vara farliga.
		-- Hawkwind

%
Det är mycket svårt att sia, särskilt när det hänför sig till framtiden.
		-- Hawkwind

%
Det är inte lätt att vara en fredag ​​typ av person i en måndag sorts värld.
		-- Hawkwind

%
Det ser ut som blinda skrikande hedonism vann.
		-- Hawkwind

%
Det slog mig nyligen att ingenting har inträffat till mig nyligen.
		-- Hawkwind

%
"Det var en urskog, en plats där Hand of Man hade aldrig satt sin fot."
		-- Hawkwind

%
Det var en av de perfekta sommardagar - solen skiner, en vindblåste, fåglarna sjunger, och gräsklipparen var bruten ...
		-- James Dent

%
Det var trevligt för mig att få ett brev från dig häromdagen. KanskeJag borde ha funnit det trevligare om jag hade kunnat tolka det. jagtror inte att jag behärskar något utöver det datum (som jag visste) ochsignaturen (som jag gissade på). Det finns en unik och en ständigcharm i ett brev till dig; det aldrig blir gammal, aldrig förlorar sinnyhet. Andra bokstäver läses och kastas bort och glömt, mendin hålls alltid - olästa. En av dem kommer att pågå en rimligmänniskan en livstid.
		-- Thomas Aldrich

%
Det var inte att hon hade en ros i tänderna, exakt. Det var mer somrosen och tänderna var i samma glas.
		-- Thomas Aldrich

%
Det skulle spara mig en hel del tid om du bara gav upp och gick galen nu.
		-- Thomas Aldrich

%
Det kommer att bli en trevlig värld om de någonsin få den färdig.
		-- Thomas Aldrich

%
Det är en 0,88 magnum - det går igenom skolan.
		-- Danny Vermin

%
Det är fantastiskt hur mycket bättre du känner när du har gett upp hoppet.
		-- Danny Vermin

%
Det är inte fallet som dödar dig, det är landning.
		-- Danny Vermin

%
Det är ganska svårt att säga vad bringa lycka; fattigdom och rikedomhar båda misslyckats.
		-- Kim Hubbard

%
Joe syster sätter spaghetti i hennes skor!
		-- Kim Hubbard

%
Gå med i marschen att spara individualitet!
		-- Kim Hubbard

%
Bara för att allt är annorlunda betyder ingenting har förändrats.
		-- Irene Peter

%
Bara ge Alice några pennor och hon kommer att stanna upptagen i timmar.
		-- Irene Peter

%
Kilroe hic erat!
		-- Irene Peter

%
Kiss me två gånger. Jag är schizofren.
		-- Irene Peter

%
Kysser en fisk är som att röka en cykel.
		-- Irene Peter

%
Knackade, inte var du i.
		-- Opportunity

%
Vet du vad jag hatar mest? Retoriska frågor.
		-- Henry N. Camp

%
L'hasard ne favorise que l'esprit förbereda.
		-- L. Pasteur

%
La-dee-dee, la-dee-dah.
		-- L. Pasteur

%
Lake Erie dog för dina synder.
		-- L. Pasteur

%
Språket är ett virus från en annan planet.
		-- William Burroughs

%
Skrattar åt dig är som drop-sparka en sårad surrfågel.
		-- William Burroughs

%
Lemmings inte blir äldre, de bara dö.
		-- William Burroughs

%
Låt den som tar steget kom ihåg att lämna tillbaka den genom tisdag.
		-- William Burroughs

%
Låt mig uttrycka det så här: i dag kommer att bli en lärande upplevelse.
		-- William Burroughs

%
Låt andra beröm antiken; Jag är glad att jag föddes i dessa.
		-- Ovid (43 B.C. - A.D. 18)

%
Låt oss påminna oss själva om att förra årets ny idé är dagens kliché.
		-- Austen Briggs

%
Liv - Älska den eller lämna den.
		-- Austen Briggs

%
Livet är vad det är, en drömmar om hämnd.
		-- Paul Gauguin

%
Livet är både svårt och tidskrävande.
		-- Paul Gauguin

%
Livet är förenat med möjligheter att hålla käften.
		-- Paul Gauguin

%
Livet är bara en skål med körsbär, men varför jag alltid få gropar?
		-- Paul Gauguin

%
Livet är som en liknelse.
		-- Paul Gauguin

%
Livet är som en analogi.
		-- Paul Gauguin

%
Livet är inte för alla.
		-- Paul Gauguin

%
Livet skulle vara acceptabelt, men för sina nöjen.
		-- G. B. Shaw

%
Som vinter snö på sommaren gräsmatta, är tids senaste tiden gått.
		-- G. B. Shaw

%
Nedskräpning är dum.
		-- Ronald Macdonald

%
Levande fasta, dö ung, och lämna en platt lapp av päls på motorvägen!
		-- The Squirrels' Motto (The "Hell's Angels of Nature")

%
Se upp! Bakom dig!
		-- The Squirrels' Motto (The "Hell's Angels of Nature")

%
Se! Framför våra ögon, är framtiden blir det förflutna.
		-- The Squirrels' Motto (The "Hell's Angels of Nature")

%
Lookie, Lookie, här kommer kaka ...
		-- Stephen Sondheim

%
Förlora dina körkort är bara Guds sätt att säga "booga, Booga!"
		-- Stephen Sondheim

%
Tappat intresset? Det är så illa jag har förlorat apati.
		-- Stephen Sondheim

%
Älskar havet? Jag dote på det - från stranden.
		-- Stephen Sondheim

%
Tur kan inte hålla en livstid, om du dör ung.
		-- Russell Banks

%
Madness tar sin tribut.
		-- Russell Banks

%
Man som faller i masugnen är säker på att känna överspända.
		-- Russell Banks

%
Man som faller i karet av smält optiskt glas gör spektakel av själv.
		-- Russell Banks

%
Man som sover i öl fat vakna klibbig.
		-- Russell Banks

%
Marigold: SvartsjukaMint: VirtueApelsin: Din renhet lika din skönhetOrchid: skönhet, praktPansy: TankarPeach Blossom: Jag är din fångePetunia: Din närvaro lugnar migVallmo: SleepRose, vilken färg som helst: LoveRose, djupröd: Bashful skamRose, singel, rosa: EnkelhetRose, thornless, alla: Tidig infästningRose, vitt: Jag är värd digRose, gul: Minskning av kärlek, ökningen av svartsjukaRosebud, vit: Girlhood, och ett hjärta okunniga om kärlekRosmarin: MinneSolros: HögmodTulpan, röd: Förklaring av kärlekTulpan, gul: Hopplös kärViolett, blått: TrofasthetViolett, vit: ModestyZinnia: Tankar om frånvarande vänner* En upp-och-ned blossom reverserar betydelsen.
		-- Russell Banks

%
Kan hundra tusen dvärgar invadera ditt hem sjunga ostliknande lounge-ödlaversioner av låtar från Trollkarlen från Oz.
		-- Russell Banks

%
Kan en Misguided Platypus lägga sina ägg i din Jockey Shorts.
		-- Russell Banks

%
Maj lopporna av tusen kamel infest armhålorna.
		-- Russell Banks

%
Må din kamel vara så snabb som vinden.
		-- Russell Banks

%
Kan tungan fastnar på gommen med styrkan av enTusen kola.
		-- Russell Banks

%
Meester, gör du vant att köpa en anka?
		-- Russell Banks

%
Minnet bör vara utgångspunkten för närvarande.
		-- Russell Banks

%
Mene, mene, tekel, upharsen.
		-- Russell Banks

%
Metermaids äta sina ungar.
		-- Russell Banks

%
Mikrobiologi Lab: Endast Staph!
		-- Russell Banks

%
Speglar bör återspegla lite innan man kastar upp bilder.
		-- Jean Cocteau

%
Moebius strippor visa dig aldrig sin baksida.
		-- Jean Cocteau

%
Moebius gör det alltid på samma sida.
		-- Jean Cocteau

%
Måndag är ett hemskt sätt att tillbringa en sjundedel av ditt liv.
		-- Jean Cocteau

%
Mest brännande frågorna generera betydligt mer värme än ljus.
		-- Jean Cocteau

%
De flesta allmänna uttalanden är falska, inklusive denna.
		-- Alexander Dumas

%
Moder Jord är inte platt!
		-- Alexander Dumas

%
Mamma är alldeles för smart för att förstå något hon inte gillar.
		-- Arnold Bennett

%
Mount Saint Helens borde ha använt jorden kontroll.
		-- Arnold Bennett

%
Måste få nära till stan - vi slår fler människor.
		-- Arnold Bennett

%
Mitt intresse är i framtiden, eftersom jag kommer att tillbringa resten av mittliv där.
		-- Arnold Bennett

%
Oj, vad du har förändrats sedan jag har förändrats.
		-- Arnold Bennett

%
"Naomi, kön vid middagstid skatter." Jag moan.Aldrig udda eller jämnt.En man, en plan, en kanal, Panama.Fru, jag är Adam.Sitt på en potatis pan, Otis.Sitt på Otis.
		-- The Mad Palindromist

%
Aldrig vara rädd för att berätta för världen vem du är.
		-- Anonymous

%
Använd aldrig "etc." - Det gör att människor tror att det finns mer där det inte finnseller att det inte finns utrymme för att lista allt, etc.
		-- Anonymous

%
Aldrig volontär för något.
		-- Lackland

%
Nya medlemmar finns ett akut behov i samhället för förhindrande avGrymhet mot dig själv. Gäller inom.
		-- Lackland

%
Nietzsche är pietzsche, men Schiller är mördare, och Goethe är moethe.
		-- Lackland

%
Ingen fågel svävar alltför hög om han svingar med sina egna vingar.
		-- William Blake

%
No guts, ingen ära.
		-- William Blake

%
Oavsett hur cynisk du får, är det omöjligt att hålla jämna steg.
		-- William Blake

%
Oavsett hur mycket du gör du aldrig göra tillräckligt.
		-- William Blake

%
Ingen liten konst är det att sova: det är nödvändigt för detta ändamål att hållavaken hela dagen.
		-- Nietzsche

%
Ingen jak alltför smutsiga; ingen container för ihålig.
		-- Nietzsche

%
Ingen någonsin dött av ugnen rå förgiftning.
		-- Nietzsche

%
Icke-determinism är inte avsett att vara rimligt.
		-- M. J. 0'Donnell

%
Icke-sequiturs gör mig äta lampskärmar.
		-- M. J. 0'Donnell

%
Nostalgi lever livet i det förflutna körfält.
		-- M. J. 0'Donnell

%
Nostalgi är inte vad det brukade vara.
		-- M. J. 0'Donnell

%
Inte skratta, inte att klaga, inte förbanna, utan att förstå.
		-- Spinoza

%
Inget kan göras i en resa.
		-- Snider

%
Ingenting botar sömnlöshet som insikten att det är dags att stiga upp.
		-- Snider

%
Ingenting är så fast trodde som det som vi stone vet.
		-- Michel de Montaigne

%
Ingenting är så ofta oåterkalleligen missade som en daglig möjlighet.
		-- Ebner-Eschenbach

%
Inget varar för evigt.Var hittar jag ingenting?
		-- Ebner-Eschenbach

%
LÄGGA MÄRKE TILL:- Hissar kommer att vara ur ORDER I DAG -(Den närmaste fungerande hiss i byggnaden tvärs över gatan.)
		-- Ebner-Eschenbach

%
Nu finns det en våldsam film med titeln "The Croquet mord" eller "MurderMed klubbor LAGD. "
		-- Shelby Friedman, WSJ.

%
Nudister är människor som bär en knapp kostymer.
		-- Shelby Friedman, WSJ.

%
O imitatörer, du slaviskt flock!
		-- Quintus Horatius Flaccus (Horace)

%
Okej, visst.
		-- Quintus Horatius Flaccus (Horace)

%
Odets, var är din udd?
		-- George S. Kaufman

%
Oh yeah? Jo, jag minns när kön var smutsiga och luften var ren.
		-- George S. Kaufman

%
Oh, ja, jag antar att detta är bara kommer att bli en av dessa livstid.
		-- George S. Kaufman

%
Oh, wow! Titta på månen!
		-- George S. Kaufman

%
När jag slutligen räknat ut alla livets svar, ändrade de frågorna.
		-- George S. Kaufman

%
Vidare genom dimman.
		-- George S. Kaufman

%
Operatör, vänligen spåra denna uppmaning och berätta var jag är.
		-- George S. Kaufman

%
Våra krukväxter har en bra känsla för humous.
		-- George S. Kaufman

%
Våra problem är så allvarliga att det bästa sättet att tala om dem ärlightheartedly.
		-- George S. Kaufman

%
Under årens lopp har jag utvecklat min känsla av deja vu så akut att nuJag kan komma ihåg saker som har * * hänt tidigare ...
		-- George S. Kaufman

%
Paranoid Club möte på fredag. Nu ... bara försöka ta reda på var!
		-- George S. Kaufman

%
Ursäkta mig medan jag skrattar.
		-- George S. Kaufman

%
Paul Revere var en tattle-tale.
		-- George S. Kaufman

%
Frid vare över detta hus, och alla som bor i den.
		-- George S. Kaufman

%
Telefonsamtal för chucky Puh.
		-- George S. Kaufman

%
Lätt som en plätt!
		-- G. S. Koblas

%
Plast ... Aluminium ... Detta är arvtagare av universum!Kött och blod har haft sin dag ... och den dagen är förbi!
		-- Green Lantern Comics

%
Vänligen hjälpa till att hålla världen ren: andra kanske vill använda den.
		-- Green Lantern Comics

%
Vänligen förbli lugn, det är ingen idé oss båda är hysterisk samtidigt.
		-- Green Lantern Comics

%
Predestination var dömd från början.
		-- Green Lantern Comics

%
Förutsägelse är mycket svårt, särskilt när det gäller framtiden.
		-- Niels Bohr

%
Bevara den gamla, men vet den nya.
		-- Niels Bohr

%
Framsteg kan ha varit bra en gång, men det har gått för länge.
		-- Ogden Nash

%
Framstegen var okej. Bara det gick för långt.
		-- James Thurber

%
Punning är det värsta last, och det finns ingen vice versa.
		-- James Thurber

%
Pyros av världen ... ANTÄNDA !!!
		-- James Thurber

%
QED.
		-- James Thurber

%
Kvacksalvare!Kvacksalvare !! Kvacksalvare!!
		-- James Thurber

%
Fråga: Är det bättre att följa reglerna tills de är ändrade ellerhjälpa till att snabba förändringen genom att bryta dem?
		-- James Thurber

%
Snabbt!! Agera som om ingenting har hänt!
		-- James Thurber

%
Quod erat demonstrandum.[Så det är bevisat. För dem som undrade WTF QED medel.]
		-- James Thurber

%
Regniga dagar och automatvapen får alltid mig.
		-- James Thurber

%
Regniga dagar och måndagar får alltid mig.
		-- James Thurber

%
Verkligheten - vad ett begrepp!
		-- Robin Williams

%
Kom ihåg att det är en omvärlden att se och njuta.
		-- Hans Liepmann

%
Kom ihåg ... det ... uhh .....
		-- Hans Liepmann

%
Kom ihåg att köra defensivt! Och naturligtvis är det bästa försvaret ett bra anfall!
		-- Hans Liepmann

%
Motstå frestelsen är lättare när du tror att du kommer förmodligen fåen ny chans senare.
		-- Hans Liepmann

%
Ring runt kragen.
		-- Hans Liepmann

%
Gummiband har galleriets ändelser!
		-- Hans Liepmann

%
Säkerhet tredje.
		-- Hans Liepmann

%
Sjömän i fartyg, segla på! Även när vi dog, andra red ut stormen.
		-- Hans Liepmann

%
Sjönk himlen för leetle lockar.
		-- Hans Liepmann

%
Santa Claus tittar!
		-- Hans Liepmann

%
Tomtenissarna är bara en massa bisatser.
		-- Hans Liepmann

%
Satir inte ser ganska på en gravsten.
		-- Hans Liepmann

%
Spara balarna!
		-- Hans Liepmann

%
Räddning valen - Harpoon en Honda.
		-- Hans Liepmann

%
Rädda valarna. Samla hela uppsättningen.
		-- Hans Liepmann

%
Se dessa två pingviner gick in i en bar, som var riktigt dum, förden andra skulle ha sett det.
		-- Hans Liepmann

%
Hon har en väckarklocka och en telefon som inte ring - de applåderar.
		-- Hans Liepmann

%
Hon är verkligen falska.
		-- Hans Liepmann

%
"Sheriff, vi måste fånga Black Bart.""Oh, ja? Vad är han ut?""Ja, han wearin en pappershatt, en pappers skjorta, pappers byxor ochpappers stövlar. ""Vad han ville ha för?""Prasslande."
		-- Hans Liepmann

%
Shirley MacLaine dog i dag i en onormal psykisk kollision idag. två freaksi en skåpbil [Åh nej !! Det är upphovsrätts polisen !!] Hennes aura-förkolnade kroppsom att vila efter ett lovtal av Jackie Collins, kollega i SAFE [Societyav asinine Flake Underhållare]. Utdrag från några av hans mer quotablekommentarer:"Verkligen en kvinna i tiden. Dessa tider, dessa tider ...""A Renaissance kvinna. Varför i 1432 ...""En man för alla årstider. Verkligen ..."Efter ceremonin, Shirley tackade hennes sörjande och förklarade hur förtjusandedet var att "få ihop" igen, förmodligen med hänvisning till att ha henne nu dödkropp gå med henne länge döda hjärna.
		-- Hans Liepmann

%
Sight är en fakultet; ser är en konst.
		-- Hans Liepmann

%
Tystnad är det element där stora saker mode sig.
		-- Thomas Carlyle

%
Tystnad är den enda kraft som finns kvar.
		-- Thomas Carlyle

%
Slang är språk som tar bort pälsen, spottar på sina händer, och går till jobbet.
		-- Thomas Carlyle

%
Sömn är för svag och sjuklig.
		-- Thomas Carlyle

%
Stryk vägen med en löpare !!
		-- Thomas Carlyle

%
Solipsists av världen ... du redan förenas.
		-- Kayvan Sylvan

%
Vissa förändringar är så långsam, du inte märker dem. Andra är så snabb,de inte märke till dig.
		-- Kayvan Sylvan

%
Vissa delar av det förflutna måste bevaras, och en del av framtiden förhindrastill varje pris.
		-- Kayvan Sylvan

%
Vissa människor lever livet i omkörningsfilen. Du är i mötande trafik.
		-- Kayvan Sylvan

%
Someday kommer vi att titta tillbaka på detta ögonblick och plöja in i en parkerad bil.
		-- Evan Davis

%
En dag får du din stora chans - eller har du redan det?
		-- Evan Davis

%
En dag, Weederman, kommer vi att titta tillbaka på allt detta och skratta ... Det kommerförmodligen en av de djupa, kusliga de som sakta bygger på enblod-ystning maniskt skrik ... men fortfarande kommer det att vara ett skratt.
		-- Mister Boffo

%
På något sätt jag nådde överskott utan att någonsin märker när jag passerartillfredsställelse.
		-- Ashleigh Brilliant

%
På något sätt, världen alltid påverkar dig mer än du påverka det.
		-- Ashleigh Brilliant

%
Ibland, är för lång för lång.
		-- Joe Crowe

%
Någonstans är något otroligt väntar på att bli känd.
		-- Carl Sagan

%
Förr eller senare måste du betala för dina synder.(De som redan har betalat kan bortse från den här cookien).
		-- Carl Sagan

%
Förlåt. Jag har glömt vad jag skulle säga.
		-- Carl Sagan

%
Förlåt. Bra försök.
		-- Carl Sagan

%
Stabilitet i sig är inget annat än en trögare rörelse.
		-- Carl Sagan

%
Stämpla ut filateli.
		-- Carl Sagan

%
Stående på huvudet gör leende rynka pannan, men resten av ansiktet också upp och ned.
		-- Carl Sagan

%
Att stjäla en noshörning bör inte försöka lätt.
		-- Carl Sagan

%
Stoppa mig, innan jag dödar igen!
		-- Carl Sagan

%
Stötta flickscouter!(Dagens Brownie är morgondagens Cookie!)
		-- Carl Sagan

%
Ta det lugnt, vi har bråttom.
		-- Carl Sagan

%
Ta vad du kan använda och låt resten gå förbi.
		-- Ken Kesey

%
Fresta mig med en sked!
		-- Ken Kesey

%
Tack för att observera alla säkerhetsföreskrifter.
		-- Ken Kesey

%
Det är konstigt. Det är mycket märkligt. Skulle inte du säga att det är mycket märkligt?
		-- Ken Kesey

%
Det är vad hon sa.
		-- Ken Kesey

%
Adjektivet är bananskal av de delar av tal.
		-- Clifton Fadiman

%
Det fina med en ordlek är i "Oy!" av betraktare.
		-- Clifton Fadiman

%
Det bästa profet framtiden är det förflutna.
		-- Clifton Fadiman

%
Vagnen har ingen plats där ett femte hjul skulle kunna användas.
		-- Herbert von Fritzlar

%
Dagen avancerade som om att tända en del arbete av mina; det var morgon,och lo! nu är det kväll, och ingenting minnesvärd uppnås.
		-- H. D. Thoreau

%
I övermorgon är den tredje dagen av resten av ditt liv.
		-- H. D. Thoreau

%
Skillnaden mellan denna plats och yoghurt är att yoghurt har ett levande kultur.
		-- H. D. Thoreau

%
Örnen kan sväva, men vesslan aldrig sugs in i en jetmotor.
		-- H. D. Thoreau

%
Bödeln är, jag hör, mycket expert, och nacken är mycket smal.
		-- Anne Boleyn

%
Det faktum att det fungerar är oväsentlig.
		-- L. Ogborn

%
... Felet som gör perfektion perfekt.
		-- L. Ogborn

%
Framtiden är inte vad den brukade vara. (Det var aldrig.)
		-- L. Ogborn

%
Framtiden ligger framför.
		-- L. Ogborn

%
Framtiden inte att födas, min vän, kommer vi att avstå från att döpa den.
		-- George Meredith

%
Gräset är alltid grönare på andra sidan av dina solglasögon.
		-- George Meredith

%
Groundhog är som de flesta andra profeter; Det levererar sitt budskap och sedanförsvinner.
		-- George Meredith

%
Förhandlingen örat finns alltid nära till den talande tunga, en anpassadvarav minnet av människan inte flöda howsomever motsatsen, SI OCH SÅ.
		-- George Meredith

%
Det viktiga att komma ihåg om att gå på ägg är inte att hoppa.
		-- George Meredith

%
"Jiggen är slut, Elman.""Vilken jigg?"
		-- Jeff Elman

%
Killer Ducks kommer !!!
		-- Jeff Elman

%
Den sista personen som sade att (Gud vila sin själ) levde att ångra det.
		-- Jeff Elman

%
Den tur som är instiftat för du kommer att bli eftertraktade av andra.
		-- Jeff Elman

%
De kanaler på mars var klart Mars sista desperat försök!
		-- Jeff Elman

%
Mygga finns att hålla den mäktiga ödmjuk.
		-- Jeff Elman

%
De viktigaste sakerna måste varje person göra för sig själv.
		-- Jeff Elman

%
En bra sak om att upprepa dina misstag är att du vet när du skakrypa.
		-- Jeff Elman

%
Det förflutna ser alltid bättre än det var. Det är bara trevligt eftersomDet är inte här.
		-- Finley Peter Dunne (Mr. Dooley)

%
Filosofen behandling av en fråga är som behandling av en sjukdom.
		-- Wittgenstein.

%
Föroreningarna är på det konstigt arrangerar. För tjock för att navigera och förtunn för att kultivera.
		-- Doug Sneyd

%
Problemet med någon oskriven lag är att du inte vet var du ska gåför att radera det.
		-- Glaser and Way

%
Läsaren meddelandet möter inte underlåta att förstå är förbannad.
		-- Glaser and Way

%
Rosen av fordom är bara ett namn, är bara namn kvar till oss.
		-- Glaser and Way

%
Fåren dog i ullen.
		-- Glaser and Way

%
Fåren som flyger över huvudet är snart att landa.
		-- Glaser and Way

%
Det kortaste avståndet mellan två godtyckliga puns är en rät linje.
		-- Glaser and Way

%
Den sjätte schejk sjätte sheeps sjuk.[Så säger den mening sextuply ...]
		-- Glaser and Way

%
Himlen är blå så vi vet var de ska sluta klippning.
		-- Judge Harold T. Stone

%
Trädet där saven är stillastående förblir fruktlös.
		-- Hosea Ballou

%
Hela jorden är i fängelse och vi rita denna fantastiska jailbreak.
		-- Wavy Gravy

%
Hela världen är en sårskorpa. Poängen är att plocka ett konstruktivt sätt.
		-- Peter Beard

%
Världen är verkligen inte något värre. Det är bara det att nyhetsbevakningenär så mycket bättre.
		-- Peter Beard

%
Världen vill bli lurade.
		-- Sebastian Brant

%
Den värsta delen av tapperhet är tanklöshet.
		-- Sebastian Brant

%
Sedan försiktigt röra mitt ansikte, tvekade hon för ett ögonblick som hennes otroögon hälls ut i min kärlek, glädje, smärta, tragedi, acceptans och fred."" Hej för nu ", sade hon varmt.
		-- Thea Alexander, "2150 A.D."

%
Det finns inga regler för mars. Mars är våren, typ av vanligen marsbetyder kanske, men inte satsa på det.
		-- Thea Alexander, "2150 A.D."

%
Det finns tre saker som jag alltid glömmer. Namn, ansikten - den tredje Ikan inte minnas.
		-- Italo Svevo

%
Det finns två typer av fotgängare ... snabbt och döda.
		-- Lord Thomas Rober Dewar

%
Det har skett en oroväckande ökning av antalet saker som du vetingenting om.
		-- Lord Thomas Rober Dewar

%
Det finns en naturlig Hootchy-Kootchy till en guldfisk.
		-- Walt Disney

%
Det finns alltid någon sämre än dig själv.
		-- Walt Disney

%
Det finns alltid något nytt ut ur Afrika.
		-- Gaius Plinius Secundus

%
Det finns inget sådant som ett problem utan en present till dig i sina händer.
		-- Gaius Plinius Secundus

%
Det finns inget nytt förutom vad som glömts bort.
		-- Marie Antoinette

%
Det verkar ingen plan eftersom det är allt plan.
		-- C. S. Lewis

%
Det finns inget behov av att göra hushållsarbete - efter fyra år det inte blirvärre.
		-- C. S. Lewis

%
Det finns inget mycket mystiskt om dig, förutom attingen riktigt vet din ursprung, syfte, eller destination.
		-- C. S. Lewis

%
De fick slutligen kung Midas, hör jag. Förgylla by association.
		-- C. S. Lewis

%
De surrade bara och surrade ... surrade.
		-- C. S. Lewis

%
Tänka stort. Förorena Mississippi.
		-- C. S. Lewis

%
Tänk tuta, om du är en telepat.
		-- C. S. Lewis

%
Tänk i sidled!
		-- Ed De Bono

%
Detta är inte en upprepning.
		-- Ed De Bono

%
Detta är i morgon du orolig igår. Och nu vet du varför.
		-- Ed De Bono

%
Detta måste vara på morgonen. Jag kunde aldrig få kläm på morgnarna.
		-- Ed De Bono

%
Denna mening motsäger sig själv - ingen faktiskt inte.
		-- Douglas Hofstadter

%
Denna mening faktiskt inte har egenskapen den påstår inte att ha.
		-- Douglas Hofstadter

%
Denna mening ingen verb.
		-- Douglas Hofstadter

%
Tre minuters trodde skulle räcka till för att ta reda på detta, men tanken ärbesvärliga och tre minuter är en lång tid.
		-- A. E. Houseman

%
Klockan tre på eftermiddagen är alltid bara en lite för sent eller liteför tidigt för allt du vill göra.
		-- Jean-Paul Sartre

%
Tid är men strömmen jag gå fiske i.
		-- Henry David Thoreau

%
Tiden kommer att avsluta alla mina bekymmer, men jag vet inte alltid godkänner Time metoder.
		-- Henry David Thoreau

%
Tis mans perdition att vara säker, när för sanningen måste han dö.
		-- Henry David Thoreau

%
Att generalisera är att vara en idiot.
		-- William Blake

%
Att älska är bra, älskar att vara svårt.
		-- William Blake

%
Att se dig är att sympatisera.
		-- William Blake

%
"Att vackla eller inte vackla, det är frågan ... eller är det?"
		-- William Blake

%
Topologists är bara plana folk.Piloter är bara plana folk.Snickare är bara plana folk.Midwest bönder är helt enkelt folk.Musiker är bara blåst folk.Deckare läsare är bara Spillane folk.Vissa Londonbor är bara P. Lane folk.
		-- William Blake

%
Problem kommer alltid vid fel tidpunkt.
		-- William Blake

%
Trouble slår i serie av tre, men när man arbetar runt husetnästa jobb efter en serie av tre är inte den fjärde jobbet - det är i början aven helt ny serie av tre.
		-- William Blake

%
Trogen vårt förflutna vi arbetar med en ärftlig, observerades och accepterade visionpersonlig fåfänga, och skönheten i världen.
		-- David Mamet

%
Två bilar i varje pott och en kyckling i varje garage.
		-- David Mamet

%
Använd en vits, gå till fängelse.
		-- David Mamet

%
Vänta för den visaste av alla rådgivare, Time.
		-- Pericles

%
Vill du köpa en anka?
		-- Pericles

%
Slösa tid är en viktig del av livet.
		-- Pericles

%
Vi har öron, Earther ... fyra av dem!
		-- Pericles

%
Vi har pågått tillräckligt länge på stranden av den kosmiska oceanen.
		-- Carl Sagan

%
Vi måste dö eftersom vi har känt dem.
		-- Ptah-hotep, 2000 B.C.

%
Vi kommer att passera den bron när vi kommer tillbaka till det senare.
		-- Ptah-hotep, 2000 B.C.

%
Välkommen till djurparken!
		-- Ptah-hotep, 2000 B.C.

%
Väl thaaaaaaat är okej.
		-- Ptah-hotep, 2000 B.C.

%
Tja, är det handskrift på golvet.
		-- Joe E. Lewis

%
Tja, vi verkligen ha en fest, men vi har gotta post en vakt utanför.
		-- Eddie Cochran, "Come On Everybody"

%
Vad som orsakar den mystiska död alla?
		-- Eddie Cochran, "Come On Everybody"

%
Vilken färg är en kameleont på en spegel?
		-- Eddie Cochran, "Come On Everybody"

%
"Vad gjorde du när skeppet sjönk?""Jag tog en kaka av tvål och tvättade mig i land."
		-- Eddie Cochran, "Come On Everybody"

%
Vad betyder "det" betyder i meningen "Vad är klockan?"?
		-- Eddie Cochran, "Come On Everybody"

%
Vad ursäkter stå i vägen? Hur kan du eliminera dem?
		-- Roger von Oech

%
Vad händer när du skära djungeln? Det avtar.
		-- Roger von Oech

%
Vad är ljudet av en hand klappar?
		-- Roger von Oech

%
Vad som snart blir gammal? Tacksamhet.
		-- Aristotle

%
	"Vad är klockan?""Jag vet inte, det håller på att förändras."
		-- Aristotle

%
Vad vi inte kan tala om vi måste passera över i tystnad.
		-- Wittgenstein

%
Vad ska du göra om alla dina problem inte löses genom den tid du dö?
		-- Wittgenstein

%
Vad du vill, vad du hänger runt i världen väntar på, är förnågot att ske till dig.[Citerat i "VMS interna och datastrukturer", V4.4, närhänvisning till AST: s.]
		-- Robert Frost

%
Vad!? Mig orolig?
		-- Alfred E. Newman

%
Vad är det här brouhaha?
		-- Alfred E. Newman

%
Vad är det som är så kul?
		-- Alfred E. Newman

%
"Vad är det för användning av en bra offert om du inte kan ändra det?"
		-- The Doctor

%
Vad hände med evig sanning?
		-- The Doctor

%
När en kamel flugor, skrattar ingen om det inte blir mycket långt!
		-- The Doctor

%
När en ko skrattar, inte mjölk kommer ut ur nosen?
		-- The Doctor

%
När en fluga landar på taket, gör den en halv rulle eller en halv loop?
		-- The Doctor

%
När blir senare blir aldrig?
		-- The Doctor

%
När man äter en elefant tar en tugga i taget.
		-- Gen. C. Abrams

%
När nöje kvarstår betyder förbli ett nöje?
		-- Gen. C. Abrams

%
När det engelska språket får i mitt sätt, jag går över den.
		-- Billy Sunday

%
När det går bra, förvänta sig något att explodera, erodera, kollaps ellerbara försvinna.
		-- Billy Sunday

%
När du slår fel nummer du aldrig få en upptagetton.
		-- Billy Sunday

%
När du är down and out, häv upp din röst och skrika, "jag ner och ut"!
		-- Billy Sunday

%
När du är redo att ge upp kampen, som kan du överlämnande till?
		-- Billy Sunday

%
När minnet går, glöm det!
		-- Billy Sunday

%
Var är jag? Vem är jag? Är jag? jag
		-- Billy Sunday

%
Var kommer det sluta? Förmodligen någonstans i närheten av där det hela började.
		-- Billy Sunday

%
Varav en inte kan tala, detta måste man vara tyst.
		-- Wittgenstein

%
Vilket är värre: okunnighet eller apati? Vem vet? Vem bryr sig?
		-- Wittgenstein

%
Piska, piska det bra!
		-- Wittgenstein

%
Vem är du?
		-- Wittgenstein

%
Vem dat som säger "vem dat" när jag säger "vem dat"?
		-- Hattie McDaniel

%
Som trasslat med min anti-paranoia skjuten?
		-- Hattie McDaniel

%
Vem kommer att ta hand om i världen när du är borta?
		-- Hattie McDaniel

%
Varför är du så svårt att ignorera?
		-- Hattie McDaniel

%
Varför måsar bor nära havet? För om de levde nära bukten,de skulle kallas baygulls.
		-- Hattie McDaniel

%
Varför ett fartyg bär last och en lastbil bära transporter?
		-- Hattie McDaniel

%
Varför kallas det en rolig ben när det gör så ont?
		-- Hattie McDaniel

%
Varför tar det så lång tid för henne att få ut allt det goda i dig?
		-- Hattie McDaniel

%
Varför finns det inte ett särskilt namn för toppar i fötterna?
		-- Lily Tomlin

%
Varför inte gå ut på en lem? Är inte det där frukten är?
		-- Lily Tomlin

%
Varför skulle någon vilja att kallas "senare"?
		-- Lily Tomlin

%
Utan äventyr, är civilisation i hela förfall.
		-- Alfred North Whitehead

%
Skulle att min hand var så snabb som min tunga.
		-- Alfieri

%
Skulle du vilja driva planlöst i min riktning?
		-- Alfieri

%
Skulle du vilja se ruinerna av mina goda avsikter?
		-- Alfieri

%
FEL!
		-- Alfieri

%
Du auto köp nu.
		-- Alfieri

%
Du kan bur en svala, kan inte du,men du kan inte svälja en bur, kan du?Flicka, bad på Bikini, kollat ​​pojke,finner pojke kollat ​​bikini på bad flicka.En man, en plan, en kanal - Panama!
		-- The Palindromist

%
Du kan komma dit härifrån, men varför i hela friden skulle du vilja?
		-- The Palindromist

%
"Du måste tänka på i morgon!""I morgon! Jag har inte ens förberett för * _________ igår * ännu!"
		-- The Palindromist

%
Zeus gav Leda fågeln.
		-- The Palindromist

%
Jo, jag tror att vi ska få några tegelstenar och vissa fladdermöss, och visa honomden * verkliga * innebörden av julen!
		-- Bernice, "Designing Women", 12/2/91.

%
Jag brukade ha mardrömmar som Grinchen hund skulle kidnappa mig och gör migklä upp i en grimma-top och hotpants och lyssna på Burl Ives poster.
		-- Robin, "Anything But Love", 12/18/91.

%
[] Skydda detta meddelande - det är en viktig historisk dokument.[] Stryk efter att ha läst - Subversive litteratur.[] Ignorera och gå tillbaka till vad du gjorde.
		-- Robin, "Anything But Love", 12/18/91.

%
Crito, jag är skyldig en kuk till Asklepios, kommer du ihåg att betala skulden?
		-- Socrates' last words

%
Jag är trött på att slåss ... De gamla män är alla döda ... De små barnfryser ihjäl. Mitt folk, en del av dem, har rymt tillkullar och har inga filtar, ingen mat. Ingen vet var de är ... Hörmig mina chefer !! Jag är trött: mitt hjärta är sjuk och ledsen. Varifrån solenNu står jag kommer att kämpa mer. Chief Joseph (Nez Perce)
		-- Socrates' last words

%
[I] f du försöker välja mellan två teorier och en ger dig enursäkt för att vara lat, är nog rätt den andra. "
		-- Paul Graham, "What You'll Wish You'd Known"

%
Oavsett om dina omslag stjärna en manlig eller en kvinnlig, jag läser din tidning förartiklar
		-- Leo Costales, in "Outside July 2005"

%
