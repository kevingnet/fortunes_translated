En Thaum är den grundläggande enheten i magiska styrka. Det har varit allmäntetablerad som den mängd av magi som behövs för att skapa en liten vit duvaeller tre normalstora biljardbollar.
		-- Terry Pratchett, "The Light Fantastic"

%
"En guide kan inte göra allt, ett faktum de flesta magiker är ovilliga att erkänna,tala diskutera med potentiella kunder. Ändå kvarstår det faktum attdet finns vissa föremål och människor, som är, för en eller annan anledning,helt immun mot någon direkt magisk trollformel. Det är för denna grupp avvarelser som magikern lär subtiliteter att använda indirekta stavar.Det gör inte heller någon skada, i att hantera dessa frågor, för att utföra en stor klubbnära din person hela tiden. "
		-- The Teachings of Ebenezum, Volume VIII

%
En forntida ordspråk sammanfattade det: när en trollkarl är trött på att leta efterkrossat glas i sin middag, det sprang, han är trött på livet.
		-- Terry Pratchett, "The Light Fantastic"

%
Kaos är kung och Magic är lös i världen.
		-- Terry Pratchett, "The Light Fantastic"

%
Rota i inte i angelägenheterna av trollkarlar, för de blir blöta och svårljus.
		-- Terry Pratchett, "The Light Fantastic"

%
Kasta inte fimpar i urinoaren, ty de är subtila ochsnar till vrede.
		-- Terry Pratchett, "The Light Fantastic"

%
"Rota i inte i angelägenheterna av guider, för du är krispigt och bramed ketchup. "
		-- Terry Pratchett, "The Light Fantastic"

%
Gör vad du vill skall vara hela lagen.
		-- Aleister Crowley

%
Åtta var även antalet Bel-Shamharoth, vilket var anledningen till en förnuftig guidenskulle aldrig nämna numret om han kunde undvika det. Eller du kommer att bli åttalevande, lärlingar skämt varnade. Bel-Shamharoth var särskiltattraherad dabblers i magi som genom att vara så det var beachcombers påstranden av onaturliga, redan halv-insnärjd i sina nät.Rincewind rumsnummer i sin inkvartering varit 7a. Han hade intevarit förvånad.
		-- Terry Pratchett, "The Sending of Eight"

%
"Hur vet du att hon är en enhörning?" Molly krävde. "Och varför var du räddatt låta henne röra dig? Jag såg dig. Du var rädd för henne. ""Jag tvivlar på att jag kommer att kännas som att prata för mycket länge," kattensvarade utan agg. "Jag skulle inte slösa tid på dårskap om jag vardu. När det gäller den första frågan, kan ingen katt ur sin första päls någonsin varalurad av framträdanden. Till skillnad från människor, som tycker om dem. Vad gäller dinandra frågan - "Här är han vacklade, och plötsligt blev mycket intresseradvid tvätt; inte heller skulle han tala förrän han slickade sig fluffig och sedanslickade sig släta igen. Även då han inte skulle titta på Molly, mensökte klorna."Om hon hade rört vid mig", sade han mycket tyst, "Jag skulle ha varithennes och inte min egen, aldrig igen. "
		-- Peter S. Beagle, "The Last Unicorn"

%
Det är ett välkänt faktum att krigare och trollkarlar inte komma överens, eftersomen sida anser den andra sidan att vara en samling av blodtörstiga idiotersom inte kan gå och tänka på samma gång, medan den andra sidan är naturligtvismisstänksamma mot en kropp av män som mumlar en hel del och bär långa klänningar. Åh, sägguiderna, om vi ska vara så, då, hur alladubbade kragar och oljade muskler Nere vid Unga Män s Pagan Association?Till vilken hjältarna svara, det är en ganska bra påstående från ett gängwimpsoes som inte kommer att gå i närheten av en kvinna på grund, kan du tro det, av derasmystisk kraft som slags dräneras ut. Höger, säger guiderna, som baraom gör det, du och din läder poserar påsar. Oh ja, säger denhjältar, varför inte du ...
		-- Terry Pratchett, "The Light Fantastic"

%
Det är väl känt att * saker * från oönskade universum söker alltiden ingång till denna, vilket är den psykiska motsvarigheten till hands förbussar och närmare till butikerna.
		-- Terry Pratchett, "The Light Fantastic"

%
Det verkar som det är det här trollkarl arbetar en av de lyxiga kryssningsfartygför ett par år. Han behöver inte ändra sina rutiner mycket som publikenförändras över ganska ofta, och han har ett bra liv. Det enda problemet ärfartygets papegoja, som sittpinnar i hallen och klockor honom natt efter natt, årefter år. Slutligen listar ut papegojan hur nästan varje trick fungerar ochbörjar ge bort för publiken. Till exempel, när magikern gören bukett blommor försvinner, papegoja squawks "bakom ryggen! Bakomryggen! "Tja, är magikern verkligen irriterad på detta, men det finns inte myckethan kan göra åt det som papegojan är en fartygs maskot och mycket populär medpassagerare.En natt, slår fartyget vissa flytande skräp, och sjunker utanett spår. Nästan alla ombord var förlorad, med undantag för magikern ochpapegoja. För tre dagar och nätter de bara driver, med magikern klängandetill en ände av en bit drivved och papegoja ligger högst upp på den andra änden.När solen går upp på morgonen den fjärde dagen, går papegojan över tillmagikerns slutet av loggen. Med uppenbara avsky i rösten, snaps han"OK, du vinner, jag ger upp. Var har du dölja skeppet?"
		-- Terry Pratchett, "The Light Fantastic"

%
Kunskap är makt - kunskap delas är energiförlust.
		-- Aleister Crowley

%
Magi är alltid den bästa lösningen - särskilt tillförlitlig magi.
		-- Aleister Crowley

%
Oavsett hur subtil guiden en kniv i skulderbladen kommer att allvarligtkramp hans stil.
		-- Aleister Crowley

%
Rincewind hade allmänt ansetts av sina lärare att vara en naturlig trollkarlpå samma sätt som fisk är naturliga bergsklättrare. Han förmodligen skulle hakastats ut ur Unseen University ändå - han kunde inte komma ihåg trollformler ochrökning gjorde honom att känna sig sjuk.
		-- Terry Pratchett, "The Light Fantastic"

%
Någonstans, precis utom synhåll, är enhörningar samla.
		-- Terry Pratchett, "The Light Fantastic"

%
Standard magiska ordet "Abracadabra", i själva verket är en förvrängning avHebreiska frasen "ha-Bracha dab'ra" som betyder "uttala välsignelsen".
		-- Terry Pratchett, "The Light Fantastic"

%
"Den första regeln av magi är enkel. Slösa inte din tid vinkahänder och hoppas när en sten eller en klubb kommer att göra. "
		-- McCloctnik the Lucid

%
De sju ögon Ningauble guiden flöt tillbaka till sin huva som hanrapporteras till Fafhrd: "Jag har sett mycket, men kan inte förklara alla The Gray.Mouser är exakt tjugofem fot under den djupaste källare i palatsetav Gilpkerio Kistomerces. Även om tjugofyra delar i tjugofemhonom är död, han lever."Nu om Lankhmar. Hon har invaderat hennes väggar brutitallt och desperat slåss pågår på gatorna, med en hårdvärd som ut-tal Lankhamar invånare från femtio till - ochutrustade med alla moderna vapen. Ändå kan du rädda staden. "	"Hur?" krävde Fafhrd.Ningauble ryckte på axlarna. "Du är en hjälte. Du bör känna till."
		-- Fritz Leiber, "The Swords of Lankhmar"

%
"Men vad är magi för?" Prince Lir krävde vilt. "Vilken nytta ärtrolldom om det inte kan spara en enhörning? "Han grep trollkarl axelhårt, för att inte falla.Schmendrick inte vända på huvudet. Med en touch av sorg hån ihans röst, sade han, "Det är vad hjältar är för."..."Ja, naturligtvis", säger han [Prince Lir] sa. "Det är precis vad hjältarär för. Wizards gör ingen skillnad, så de säger att ingenting gör, menhjältar är avsedda att dö för enhörningar. "
		-- Peter Beagle, "The Last Unicorn"

%
Det finns de som hävdar att magi är som tidvattnet; att den sväller ochbleknar över jordens yta, samla i koncentrerade pooler häroch där, nästan försvinner från andra platser, lämnar dem torra förundra. Det finns också de som tror att om du håller fingrarna uppnäsan och blåsa, kommer det att öka din intelligens.
		-- The Teachings of Ebenezum, Volume VII

%
Unseen University hade aldrig erkänt kvinnor, muttrade något omproblem med VVS, men det verkliga skälet var en outtalad fruktan somom kvinnor tilläts röra runt med magi skulle de förmodligen varapinsamt bra på det ...
		-- Terry Pratchett, "The Light Fantastic"

%
Använda ord för att beskriva magi är som att använda en skruvmejsel för att skära rostbiff.
		-- Tom Robbins

%
"Sannerligen och forsooth", svarade Goodgulf mörkt. "Under det senaste åretkonstiga och rädda undrar jag har sett. Fält sådda med korn skördacrabgrass och svamp, och även små trädgårdar avvisar deras kronärtskocka hjärtan.Det har varit en varm dag i december och en blå måne. Kalendrar är gjorda meden månad av söndagar och en blå-band Holstein bar levande två försäkringförsäljare. Jorden splittringar och inälvorna av en get hittades bunden ikvadratiska knop. Inför solen svartnar och himlen har regnat nerfuktig chips. ""Men vad gör alla dessa saker detta?" flämtade Frito."Slår mig", sa Goodgulf med en axelryckning, "men jag tyckte det gjorde brakopiera."
		-- Harvard Lampoon, "Bored of the Rings"

%
Titta Rincewind.Titta på honom. Magra, liksom de flesta guider, och klädd i en mörkröd mantel påsom några mystiska sigils var broderade i skamfilat paljetter. vissa kanskehar tagit honom för en enkel lärling trollkarl som hade rymt från sinmästare av trots, tristess, rädsla och en kvardröjande smak förheterosexualitet. Ändå runt halsen var en kedja som bär brons oktagonsom markerade honom som en före detta elev av osedda universitet, high school av magivars tid och rymd transcendenta campus är aldrig exakt här eller där.Examinerade var oftast avsett för mageship minst, men Rincewind - efteren olycklig händelse - hade lämnat veta endast en stava och gjorde en levande avsorterar runt staden genom att utnyttja en medfödd gåva för språk. hanundvek arbete som regel, men hade en snabbhet av intelligens som lade sinbekanta i huvudet på en ljus gnagare.
		-- Terry Pratchett, "The Colour of Magic"

%
Vad är en trollkarl, men en praktiserande teoretiker?
		-- Obi-Wan Kenobi

%
Vilken nytta är magiskt om det inte kan spara en enhörning?
		-- Peter S. Beagle, "The Last Unicorn"

%
När jag säger det magiska ordet till alla dessa människor, kommer de att försvinna för alltid.Jag kommer då att säga de magiska orden för dig, och du kommer också att försvinna - aldrigses igen.
		-- Kurt Vonnegut Jr., "Between Time and Timbuktu"

%
