En karriär är stor, men du kan inte köra fingrarna genom sitt hår.
		-- Pat Benatar, "Hell is for Children"

%
En kyss är en kurs av förfarande, listigt utformas, för ömsesidigtstopp för tal vid en tidpunkt då ord är överflödiga.
		-- Pat Benatar, "Hell is for Children"

%
En kvinna var kär i fjorton soldater. Det var helt klart platoonic.
		-- Pat Benatar, "Hell is for Children"

%
Frånvaro minskar mediokra passioner och ökar stora sådana,som vinden blåser ut ljusen och fläktar bränder.
		-- La Rochefoucauld

%
Frånvaro i kärlek är som vatten på eld; lite quickens, men mycketsläcker den.
		-- Hannah More

%
Alla passioner gör oss begå fel; kärlek gör oss begå mestlöjligt sådana.
		-- La Rochefoucauld

%
Alltid kvarstår delar av vårt hjärta, i vilken ingen kan komma in,bjuda in dem som vi kan.
		-- La Rochefoucauld

%
Bondage kanske, disciplin aldrig!
		-- T.K.

%
Misstro alla dem som älskar dig mycket på en mycket liten bekantskapoch utan någon synlig orsak.
		-- Lord Chesterfield

%
Misströsta inte, din ideala älskare väntar på dig runt hörnet.
		-- Lord Chesterfield

%
Falling in LoveNär två personer har varit på tillräckligt många datum, de i allmänhet faller ikärlek. Du kan tala om du är kär i hur du känner: huvudet blirljus, hoppar ditt hjärta inom dig, du känner att du går på luft,och hela världen verkar vara en underbar och glad plats. Tyvärr,Dessa är också de fyra varningstecken kolon sjukdom, så det är alltid enbra idé att kontrollera med din läkare.
		-- Dave Barry

%
Falling in love är en mycket som dör. Du får aldrig göra det tillräckligt för attbli bra på det.
		-- Dave Barry

%
Avsluta meningen nedan i 25 ord eller mindre:"Kärlek är vad du känner precis innan du ger någon en bra ..."Post ditt svar tillsammans med den övre halvan av din handledare till:P.O. Box 35Förbryllad grekiska, Michigan
		-- Dave Barry

%
Ge mig kyskhet och continence, men inte just nu.
		-- St. Augustine

%
Gud är kärlek, men få det skriftligt.
		-- Gypsy Rose Lee

%
"Han bestämmer dock att med mer tid och en hel del mentalansträngning, kunde han förmodligen vända verksamheten till en acceptabel perversion. "
		-- Mick Farren, "When Gravity Fails"

%
Han som är kär i sig själv har åtminstone denna fördel - han kommer intemöter många konkurrenter.
		-- Georg Lichtenberg, "Aphorisms"

%
Hjärtan kommer aldrig att vara praktiska, tills de kan göras unbreakable.
		-- The Wizard of Oz

%
HEY KIDS! ANN LANDERS SÄGER:Var säker på att det är sant, när du säger "jag älskar dig". Det är synd att	berätta en lögn. Miljontals hjärtan har brutits, bara för attdessa ord uttalades.
		-- The Wizard of Oz

%
Hans hjärta var ditt från första stund som du träffade.
		-- The Wizard of Oz

%
Hur mycket hon älskar dig? Mindre än du någonsin kommer att veta.
		-- The Wizard of Oz

%
Jag är två dårar, jag vet, för att älska, och för att säga så.
		-- John Donne

%
Jag kan laga pausen på dagen, läka ett brustet hjärta, och ge tillfälligtlättnad för nymfomaner.
		-- Larry Lee

%
Jag vill inte att folk ska älska mig. Det gör för skyldigheter.
		-- Jean Anouilh

%
Jag älskar dig mer än något i denna värld. Jag tror inte att kommer att pågå.
		-- Elvis Costello

%
Jag älskar dig, inte bara för vad du är, men för vad jag är när jag är med dig.
		-- Roy Croft

%
Jag älskade henne med en kärlek törstig och desperat. Jag kände att vi två skulle begånågra agera så fruktansvärda att världen, se oss, skulle finna det oemotståndliga.
		-- Gene Wolfe, "The Shadow of the Torturer"

%
Jag har aldrig älskat en annan person som jag älskade mig.
		-- Mae West

%
Jag tror att en relation är som en haj. Det måste hela tiden gå framåteller det dör. Nå, vad vi har på våra händer här är en död haj.
		-- Woody Allen

%
Jag brukade vara Snövit, men jag drev.
		-- Mae West

%
Jag brukade tänka romantisk kärlek var en neuros som delas av två, en högstadåraktighet. Jag trodde inte längre det. Det finns inget dumtkärleksfull någon. Tänker du bli älskad i gengäld är det är dumt.
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag gjorde min egen grej och nu har jag fåttatt ångra det. "
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag måste tandtråd min katt."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag måste stanna hemma och se om jag snarkar."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag går aldrig ut på dagar som slutar på 'Y.'"
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag vill tillbringa mer tid med min mixer."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag närvara vid öppnandet av min garageport."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag omvandla min kalender klocka frånJulian till gregorianska. "
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag gör dörr till dörr insamling för statiskhålla fast."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag har alla mina växter kastrerad."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag stannar hemma för att arbeta på minkeso skulptur. "
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag tar punk totempåle carving."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men jag har planerat för en karma transplantation."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men det är min undulat bowling kväll."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men min favorit kommersiella är på tv."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men förra gången jag gick ut, aldrig kom jag tillbaka."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men mannen på TV berättade för mig att hålla ögonen öppna."
		-- Rita Mae Brown

%
"Jag skulle gärna vilja gå ut med dig, men det finns viktiga världsfrågor sombehöver oroa dig. "
		-- Rita Mae Brown

%
Jag vill gärna kyssa dig, men jag tvättade bara mitt hår.
		-- Bette Davis, "Cabin in the Cotton"

%
"Jag ska berätta vad jag vet, då," han bestämt. "Stiftet jag bärbetyder att jag är medlem i IA. Det är Inamorati Anonym. En inamorato ärnågon kär. Det är det värsta missbruk av alla. ""Någon är på väg att falla i kärlek" Oedipa sa, "du går sitta meddem, eller något? ""Just det. Hela idén är att komma dit du inte behöver det. Jag vartur. Jag sparkade det unga. Men det finns sextio-åriga män, tro det ellerinte, och kvinnor ännu äldre, som kanske vaknar på natten skriker. ""Du håller möten, då, i likhet med AA?""Nej, naturligtvis inte. Du får ett telefonnummer, en telefonsvararedu kan ringa. Ingen vet någon annans namn; bara antalet i falletdet blir så dålig att du inte kan hantera det ensam. Vi är isolat, Arnold. mötenskulle förstöra hela poängen med det. "
		-- Thomas Pynchon, "The Crying of Lot 49"

%
Om kärlek är svaret, kan du förtydliga frågan?
		-- Lily Tomlin

%
Om kärlek Var olja, skulle jag vara om en Quart Låg
		-- Book title by Lewis Grizzard

%
Om ni bara visste att hon älskade dig, kan du möta osäkerheten iom du älskar henne.
		-- Book title by Lewis Grizzard

%
Om du inte kan vara bra, vara försiktig. Om du inte kan vara försiktig, ge mig ett samtal.
		-- Book title by Lewis Grizzard

%
Om du älskar någon, befria dem.Om de inte kommer tillbaka, sedan ringa upp dem när du är full.
		-- Book title by Lewis Grizzard

%
I en stor roman, varje person spelar i princip en del attandra verkligen gillar.
		-- Elizabeth Ashley

%
I en tid när mode är att vara kär i dig själv, bekänna tillvara kär i någon annan är ett erkännande av otrohet till sinälskad.
		-- Russell Baker

%
Kär, hon som ger henne porträtt lovar originalet.
		-- Bruton

%
I verklig kärlek du vill att den andra personen är bra. I romantisk kärlek duvill att den andra personen.
		-- Margaret Anderson

%
Det är mycket bättre att luras än att undeceived av dem vi älskar.
		-- Margaret Anderson

%
Hur svårt det är att skriva biografi kan räkna med någonsom sitter ner och anser hur många vet den verkliga sanningenom hans eller hennes kärleksaffärer.
		-- Rebecca West

%
Låt oss leva !!!Låt oss älska !!!Låt oss dela djupaste hemligheter våra själar !!!Du först.
		-- Rebecca West

%
Låt oss bara vara vänner och göra någon särskild ansträngning för att någonsin se varandra igen.
		-- Rebecca West

%
Låt oss inte komplicera vår relation genom att försöka kommunicera med varandra.
		-- Rebecca West

%
Ensam är en man utan kärlek.
		-- Englebert Humperdinck

%
Kärlek - den sista av de allvarliga sjukdomar i barndomen.
		-- Englebert Humperdinck

%
Kärlek och skandal är de bästa sötningsmedel av te.
		-- Englebert Humperdinck

%
Kärlek vid första ögonkastet är en av de största arbetsbesparande anordningarvärlden någonsin har sett.
		-- Englebert Humperdinck

%
Kärlek kan inte vara mycket yngre än lusten för mord.
		-- Sigmund Freud

%
Kärleken övervinner allt saker; Låt oss också ge efter för kärleken.
		-- Publius Vergilius Maro (Virgil)

%
Kärlek är en allvarlig psykisk sjukdom.
		-- Plato

%
Kärlek är en snöskoter racing över tundran, som plötsligt vänderöver, sätter du nedanför. På natten isen vesslor komma.
		-- Matt Groening, "Love is Hell"

%
Kärlek är alltid öppna armar. Med öppna armar du tillåter älskar att komma ochgå som det vill, fritt, för det kommer att göra det ändå. Om du stängerarmarna om älskar dig hittar du kvar bara håller dig själv.
		-- Matt Groening, "Love is Hell"

%
Kärleken är dum tillsammans.
		-- Paul Valery

%
Kärlek är dope, inte kycklingsoppa. Jag menar, kärlek är något som ska skickasrunt fritt, inte sked ner någons hals för deras eget bästa med enJudisk mor som tillagas allt själv.
		-- Paul Valery

%
Kärlek är i görningen.
		-- The Homicidal Maniac

%
Kärlek är som en vänskap fattade eld. I början en flamma, mycketsöt, ofta varm och hård, men fortfarande bara ljus och flimmer. som kärlekblir äldre, våra hjärtan mogna och vår kärlek blir som kol, djupt bränningoch outsläcklig.
		-- Bruce Lee

%
Kärlek är som mässlingen; vi alla måste gå igenom det.
		-- Jerome K. Jerome

%
Kärlek är aldrig frågar varför?
		-- Jerome K. Jerome

%
Kärlek är inte tillräckligt, men det säkert hjälper.
		-- Jerome K. Jerome

%
Kärlek är sentimentala mässling.
		-- Jerome K. Jerome

%
Kärleken stanna uppe hela natten med ett sjukt barn, eller en frisk vuxen.
		-- Jerome K. Jerome

%
Kärlek är det enda spelet som inte kallas på grund av mörker.
		-- M. Hirschfield

%
Kärlek är den process av min leder dig försiktigt tillbaka till dig själv.
		-- Saint Exupery

%
Kärlek är en triumf för fantasin över intelligens.
		-- H. L. Mencken

%
Kärlek är vad det är knäckt upp vara.
		-- H. L. Mencken

%
Kärlek är vad du har gått igenom med någon.
		-- James Thurber

%
Kärlek är inte bara blind, det är också döv, stum och dum.
		-- James Thurber

%
Kärlek innebär med att säga att du är ledsen var femte minut.
		-- James Thurber

%
Kärlek innebär aldrig behöva säga att du är ledsen.Det är det löjligaste jag någonsin har hört.
		-- Ryan O'Neill, "What's Up Doc?"

%
Kärlek berättar många saker som inte är så.
		-- Krainian Proverb

%
Må din SO alltid vet när du behöver en kram.
		-- Krainian Proverb

%
"Kanske borde vi tänka på detta som en perfekt vecka ... där vi funnit varandraandra och älskade varandra ... och sedan låta varandra gå innan någonvar tvungen att söka professionell hjälp. "
		-- Krainian Proverb

%
De flesta människor behöver inte en stor kärlek nästan så mycket som de behöveren stadig leverans.
		-- Krainian Proverb

%
Min kopp hath runneth'd över med kärlek.
		-- Krainian Proverb

%
Naturen avskyr en jungfru - en fryst tillgångar.
		-- Clare Booth Luce

%
"Nej, jag förstår nu" Auberon sade, lugn i skogen - det var såenkel, verkligen. "Jag gjorde inte, under en lång tid, men jag gör nu. Du kan bara intehålla människor, kan du inte äger dem. Jag menar att det är naturligt, en naturlig processverkligen. Träffa. Kärlek. Del. Livet går vidare. Det var aldrig någon anledning attatt hon skulle stanna alltid samma - jag menar 'kär, "du vet" Det fanns.dessa tvivel-citat av Smoky, tungt anges. "Jag inte hålla ett agg. Ikan inte.""Du gör", sa farfar öring. "Och du inte förstår."
		-- Little, Big, "John Crowley"

%
Av alla former av försiktighet, är försiktighet älskar mest dödliga.
		-- Little, Big, "John Crowley"

%
Naturligtvis är det möjligt att älska en människa om du inte känner dem alltför väl.
		-- Charles Bukowski

%
Åh, är kärlek verkliga nog, du kommer att finna det en dag, men det har enärkefiende - och det är liv.
		-- Jean Anouilh, "Ardele"

%
På en tous un peu peur de l'amour, mais på en surtout peur de souffrirou de faire souffrir.[One är alltid lite rädd för kärlek, men framför allt en ärrädd för smärta eller orsaka smärta.]
		-- Jean Anouilh, "Ardele"

%
När insikten har accepterat att även mellan de närmaste människoroändliga avstånd fortsätter att existera, en underbar lever sida vid sida kanväxa upp, om de lyckas älska avståndet mellan dem, vilket gör detmöjligt för var och en se varandra hela mot himlen.
		-- Rainer Rilke

%
Man uttrycker väl den kärlek han inte känner.
		-- J. A. Karr

%
Folk tror att kärlek är en känsla. Kärlek är sunt förnuft.
		-- Ken Kesey

%
Verkligen?? Vilket sammanträffande, jag är för grunt !!
		-- Ken Kesey

%
Någon gång när du minst anar det, kommer att älska peka dig på axeln ...och ber dig att flytta ut ur vägen eftersom det fortfarande inte är din tur.
		-- N. V. Plyter

%
Ibland är kärlek inte bara ett missförstånd mellan två dårar.
		-- N. V. Plyter

%
Tyvärr aldrig innebär att ha din kommentar att älska.
		-- N. V. Plyter

%
På tal om kärlek, ett problem som återkommer allt oftare dessadagar, i böcker och pjäser och filmer, är oförmågan hos människor att kommuniceramed de människor de älskar; Män och hustrur som inte kan kommunicera, barnsom inte kan kommunicera med sina föräldrar, och så vidare. Och tecknen idessa böcker och pjäser och så vidare (och i verkliga livet, kan jag tillägga) tillbringar timmarbemoaning det faktum att de inte kan kommunicera. Jag tror att om en person inte kankommunicera, mycket _____ stone han kan göra är att hålla käften!
		-- Tom Lehrer, "That Was the Year that Was"

%
Support djurliv - rösta för en orgie.
		-- Tom Lehrer, "That Was the Year that Was"

%
Det är den sanna säsongen av kärlek, när vi tror att vi bara kan älska,att ingen kunde ha älskat så framför oss, och att ingen kommer att älskapå samma sätt som oss.
		-- Johann Wolfgang von Goethe

%
Det är livet för dig, sade McDunn. Någon alltid väntar på någon somaldrig kommer hem. Alltid någon kärleksfull något mer än det där älskardem. Och efter ett tag du vill förstöra vad det är, så detkan inte skada dig längre.
		-- R. Bradbury, "The Fog Horn"

%
Fåglarna sjunger, blommorna spirande, och det är dagsför Miss Manners att berätta unga älskande att sluta insnörning offentligt.Det är inte att fröken Manners är immun mot romantik. miss Mannershar varit kända för att pressa en herre arm samtidigt som hjälpt över enbromsa, och i hennes vilda ungdom, även trycka på en prydlig toffel mot enfot eller två under middagsbordet. Miss Manners anser också attåsynen av människor längsmed hand i hand eller arm i armen eller arm i handenklär upp en stad betydligt mer än de mer välkända åsynen avskakar paraplyer på varandra. Vad fröken Manners motsätter sigär den typ av aktivitet som skrämmer hästarna på gatan ...
		-- R. Bradbury, "The Fog Horn"

%
Giraffen du trodde att du kränkt förra veckan är villig att nuzzled idag.
		-- R. Bradbury, "The Fog Horn"

%
Hjärtat har sina skäl varför vet ingenting om.
		-- Blaise Pascal

%
Hjärtat är klokare än intellektet.
		-- Blaise Pascal

%
De små bitar av mitt liv jag ger till dig, med kärlek att göra ett täckeatt hålla bort kylan.
		-- Blaise Pascal

%
Det magiska av vår första kärlek är vår okunnighet som det någonsin kan sluta.
		-- Benjamin Disraeli

%
Myten om romantisk kärlek anser att när du har blivit kär i denperfekt partner, du är hemma gratis. Tyvärr faller av kärlekverkar vara lika ofrivillig falla in i den.
		-- Benjamin Disraeli

%
Den enda skillnaden i spelet av kärlek under de senaste några tusen årär att de har ändrat trumf från klubbar till diamanter.
		-- The Indianapolis Star

%
Uppkomsten och avtagande av kärlek gör sig gällande i oroerfarna vid att vara ensam tillsammans.
		-- Jean de la Bruyere

%
Den perfekta älskare är en som förvandlas till en pizza på 4:00
		-- Charles Pierce

%
Den person du avvisade igår kan göra dig lycklig, om du säger ja.
		-- Charles Pierce

%
Den sju år klådan kommer från lurar runt under fjärde, femte,och sjätte år.
		-- Charles Pierce

%
Historien om fjärilen:"Jag var i Bogota och väntar på en väninna. Jag var kär,för länge sedan. Jag väntade tre dagar. Jag var hungrig men kunde inte gåut mat, så att hon kommer och jag inte vara där för att hälsa henne. Sedan, påden tredje dagen, hörde jag en knackning. ""Jag skyndade längs den gamla kanalen och där, i solskenet,det fanns ingenting. ""Bara" Vance Joy sade, "en fjäril, flyga iväg."
		-- Peter Carey, BLISS

%
Den sötare äpplet, den svartare kärnan -Skrapa en älskare och hitta en fiende!
		-- Dorothy Parker, "Ballad of a Great Weariness"

%
Sättet att älska något är att inse att det kan gå förlorad.
		-- Dorothy Parker, "Ballad of a Great Weariness"

%
Det finns några mikroorganismer som uppvisar egenskaper hos båda anläggningarnaoch djur. När de utsätts för ljus de genomgår fotosyntes; och närljuset slocknar, de förvandlas till djur. Men återigen, inte vi alla?
		-- Dorothy Parker, "Ballad of a Great Weariness"

%
Det finns ingen rädsla i kärleken, utan fullkomlig kärlek driver ut rädsla.
		-- 1 John 4:18

%
Det finns bara ett sätt att bli lycklig genom hjärtat - att ha någon.
		-- Paul Bourget

%
Det finns så mycket att säga, men dina ögon hålla avbryter mig.
		-- Paul Bourget

%
Timing måste vara perfekt nu. Två timing måste vara bättre än perfekt.
		-- Paul Bourget

%
Att bli älskad är mycket demoraliserande.
		-- Katharine Hepburn

%
Att frukta kärlek är att frukta livet, och de som är rädda liv är redan tredelar död.
		-- Bertrand Russell

%
Totala främlingar behöver kärlek, alltför; och jag är främling än de flesta.
		-- Bertrand Russell

%
Sann lycka kommer att hittas endast i sann kärlek.
		-- Bertrand Russell

%
Under deadline tryck för nästa vecka. Om du vill ha något, kan det vänta.Om det inte är blinda skrikande paroxysmally hedonistiska ...
		-- Bertrand Russell

%
Vi tror inte på reumatism och sann kärlek förrän efter den första attacken.
		-- Marie Ebner von Eschenbach

%
Vad är irriterande om kärlek är att det är ett brott som kräver en medbrottsling.
		-- Charles Baudelaire

%
När ditt liv är ett löv som årstiderna riva av och fördömaDe kommer att binda dig med kärlek som är graciös och grönt som en stam.
		-- Leonard Cohen, "Sisters of Mercy"

%
Varför jag inte kan gå ut med dig:Jag skulle gärna vilja, men ...- Jag måste tandtråd min katt.- Jag har vigt mitt liv åt linguini.- Jag behöver spendera mer tid med min mixer.- Det skulle inte vara rättvist att andra Vackra människor.- Det är min natt att klappa hunden / iller / guldfisk.- Jag ska på stan för att prova på vissa handskar.- Jag måste kolla färskhet datum på min mejeriprodukter.- Jag ska ner till bageriet för att titta på bullarna stiga.- Jag har ett möte med en nagelband specialist.- Jag har några riktigt hårda ord för att leta upp.- Jag har fått en Friends of the Lowly Rutabaga mötet.
		-- I promised to help a friend fold road maps.

%
Varför jag inte kan gå ut med dig:Jag skulle gärna vilja, men ...- Jag måste svara på alla mina "åkandes" bokstäver.- Ingen av mina strumpor match.- Jag har alla mina växter kastrerade.- Jag bytte lås på min dörr och nu kan jag inte komma ut.- Min yucca anläggningen känner äckligt.- Jag turnerade Kina med en wok band.- Min choklad uppskattning klass möter den natten.- Jag kör iväg till Jugoslavien med ett utländskt utbytesstudentnamngav Basil Metabolism.- Det finns viktiga världsfrågor som behöver oroa.- Jag kommer att räkna borsten i min tandborste.- Jag föredrar att förbli en gåta.- Jag tror att du vill att de andra Peggy / Cathy / Mike / vem.
		-- I feel a song coming on.

%
Varför jag inte kan gå ut med dig:Jag skulle gärna vilja, men ...- Jag måste dra "Cubby" för en konststipendium.- Jag måste sitta upp med en sjuk ant.- Jag försöker att vara mindre populär.- Min badrumskakel behöver injektering.- Jag väntar på att se om jag redan en vinnare.- Min medvetna säger nej.- Jag plockade bara upp en bok som heter "Glue i många länder", och jagverkar inte kunna lägga ner.- Min favorit kommersiella är på TV.- Jag måste studera för mitt blodprov.- Jag har handlats till Cincinnati.- Jag har mina barn skor brons.
		-- I have to go to court for kitty littering.

%
Varför jag inte kan gå ut med dig:Jag skulle gärna vilja, men ...- Jag försöker att se hur länge jag kan gå utan att säga ja.- Jag närvara vid öppnandet av min garageport.- Monstren har inte vänt blå ännu, och jag måste äta fler punkter.- Jag konvertera min kalender klocka från Julian till gregorianska.- Jag måste uppfylla min potential.- Jag vill inte lämna min komfortzon.- Det är för nära sekelskiftet.- Jag måste bleka min hare.- Jag är orolig för min vertikala hålla ratten.
		-- I left my body in my other clothes.

%
Varför jag inte kan gå ut med dig:Jag skulle gärna vilja, men ...- Jag har fått en Friends of the Lowly Rutabaga mötet.- Jag lovade att hjälpa en vän vika vägkartor.- Jag har planerat för en karma transplantation.- Jag stannar hemma för att arbeta på min keso skulptur.- Det är min undulat bowling kväll.- Jag ska bygga en anläggning från ett kit.- Det finns en störning i Kraften.- Jag gör dörr till dörr insamling för statisk klänga.- Jag undervisar min iller att joddla.
		-- My crayons all melted together.

%
"Varför måste du berätta alla dina hemligheter när det är svårt nog att älskadu vet ingenting? "
		-- Lloyd Cole and the Commotions

%
Utan kärlek intelligens är farlig;utan intelligens kärlek är inte tillräckligt.
		-- Ashley Montagu

%
Skulle inte detta vara en stor värld om att osäkra och desperat var en turn-on?
		-- "Broadcast News"

%
Ja, det finns viktigare saker i livet än pengar, men de kommer inte att gåut med dig om du inte har någon.
		-- "Broadcast News"

%
Du ska inte behöva betala för din kärlek med dina ben och din kropp.
		-- Pat Benatar, "Hell is for Children"

%
