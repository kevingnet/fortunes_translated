Jag tycker det är lite fantastiskt att försöka bilda en bild i människorssinnen Debianarkivet administration laget kröp över derasterminaler, tände sina ansikten endast en CRT med en liten rot skalsnabb och kommandot"/project/org/ftp.debian.org/cabal/s3kr1t/nuke-non-free.pl" Alla knappati och redo att gå, deras fingrar redo över Enter, en svettvällustig förväntade beading på sina övre läppar. "<20031104211846.GK13131@deadbeast.net> diskuterarsitt förslag till sociala kontrakt ändring
		-- Branden Robinson in

%
Om du ska köra en rinky-dink distro som gjorts av ett parvolontärer, varför inte köra en rinky-dink distro som gjorts av en hel del frivilliga?
		-- Jaldhar H. Vyas on debian-devel

%
Förpackningarna ska bygga beror på vad de ska bygga beroende.
		-- Santiago Vila on debian-devel

%
Det finns 3 typer av killar - de som hatar nerds (alla nördar, attär; flickor inte låta undan); de som är rädd av flickorsom är något mer intelligent än genomsnittet; och killarna som ärockså något mer intelligent än genomsnittet, men är så blyg att dekan inte sätta 2 ord tillsammans när de är inom 20 fot av en flicka.
		-- Vikki Roemer on debian-curiosa

%
Debian är Jedi operativsystemet: "Alltid två finns en master ochen lärling ".
		-- Simon Richter on debian-devel

%
Detta är Unix vi pratar om, kom ihåg. Det är inte tänkt att varatrevligt för applikationer programmerare.
		-- Matthew Danish on debian-devel

%
... Men hey, detta är Linux, är det inte tänkt att göra oändliga loopar i 5sekunder?
		-- Jonathan Oxer in the apt-cacher ChangeLog

%
Jag är personligen ganska nöjd med en stabil utgåva vartannat år, ochär av den åsikten att försöka frigöra mer kommer att innebära att vi måstebyta namn på distro från "stabil" till "vinglig".
		-- Scott James Remnant on debian-devel

%
<Keybuk> Perl 6 skrämmer mig<Doogie> kan du namnge din operatörer någonting. namnet här är den          string "~ | _ | ~"* Lo-lan-2 flyr skrikande<Keybuk> det ser ut som ett diagram över en kanal lås :)<Jaybonci> japansk Smiley operatörer?<Nickr> ^ _ ^
		-- in #debian-devel

%
<Sam> /.ing ett problem är som att be ett oändligt antal apor för       råd
		-- in #debian-devel

%
<Daniels> fortfarande tron ​​blod låter som en film om overfiend           och oskulder eller någon skit
		-- in #debian-devel

%
<Jaybonci> faktiskt d-i står för "gudomligt ingripande";)
		-- in #debian-devel

%
<Doogie> asuffield: hur tror du dpkg skrevs ursprungligen? : |<Asuffield> genom att låta IWJ få farligt nära en dator
		-- in #debian-devel

%
<Asuffield> en arbetsstation är något du kan hålla på somebodies skrivbord             och con dem till att använda
		-- in #debian-devel

%
<Joshk> joshk @ tillströmning: /etc/logrotate.d> sh -n *<Joshk> apache: linje 14: syntaxfel nära oväntade token '}'<Joshk> apache: linje 14: `}"<Joshk> tomten tjocknar<Asuffield> de är inte skalskript<Erich> detta inte var kyckling.
		-- in #debian-devel

%
Jag attackerades av dselect som ett litet barn och har sedan undvikitdebian.
		-- Andrew Morton

%
* Joeyh installerar debian med enbart hans stortå, för en förändring av takten
		-- in #debian-boot

%
* Liiwi tar piska och ögon PASC<PASC> bonitooooo !!! kinky!<PASC> hur bekvämt, jag var bara om att kalla in sjuka på jobbet ;-)
		-- in #debian-devel

%
<Mörk> Det visade sig att grep returnerar felkod 1 när det inte finns några matcher.       Jag visste att. Varför tog det mig en halvtimme?
		-- Seen on #Debian

%
Det är helt enkelt otroligt hur mycket energi och kreativitet människor harinvesteras i att skapa motsägelsefulla, falska och dumma licenser ...
		-- - Sven Rudolph about licences in debian/non-free.

%
<Overfiend> partycle: jag på allvar behöver en semester från detta            paket. Jag hade faktiskt en dröm om att införa en            dum ny bugg i xbase-preinst går kväll. Det är en            Dåligt tecken.
		-- Seen on #Debian shortly before the release of Debian 2.0

%
<Mörk> Ser ut som kanalen är tillbaka till det normala :)<Jim> Du menar det inte rulla snabbare än någon kan läsa? :)
		-- Seen on #Debian after the release of Debian 2.0

%
Bara för att expandera på vad Ross sagt, det är utan tvekan mycket att väntavarje fördelning som det automatiskt detektera om eller inteperson som installerar den kan läsa enkla engelska riktningar, och om hankan inte fortsätta utan hans ingång. På så sätt ligger galenskap.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Zedboy> dackel: i allmänhet * bara * sättet att använda ett datorprogram         är att verkställa det. har du * någonsin * känt ett system verktyg vars         dokumentation rekommenderas antingen ta bort den, eller kasta den         på en gård djur?<Dackel> zedboy: Eeeh ... ja<Zedboy> dackel: installera manualsidor paketet. Det borde vara där         redan Tho.<Zedboy> dackel: exempel på en sådan bovint användbarhet?* Greycat vill ha en video från dackel kasta / usr / bin / fil på en ko
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Elmo> Joy: tack, glädje<Doogie> elmo: det är överflödigt, elmo<Elmo> doogie: gå spela i trafiken<Doogie> ah, elmo vi känner och älskar
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Doogie> glädje / elmo: varför kan inte samma ip användas? var denna brand så         stor att det brände IP-adress?
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Donnerjack> Ingenting säger "Jag trivs med dig" som gåva             3: e gradens brännskador ...<Mephron> utom naturligtvis vända sin säng i en Trebuchet.<Ladegard> Så mycket ansträngning måste betyda något slags tillgivenhet.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Bräcklig> Någon här kunnig i frågor som andfåglar? om du         promenad genom en park, och en gås börjar efter dig ... och         hamnar följer dig mer än en halv mil tills du når         bilen ... vid 11:00. Är gåsen rabiat eller något?
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Wolfgang> problemet med "gå hitta en riktig flicka" förmaning är           att så få av dem har faktiskt naken transformation           sekvenser<Verklighet> Dude, ändrar min flickvän som fyra gånger om dagen
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Z-Gryphon> Om Unicron hade en teknisk spec kort, skulle hans motto vara "Det            som inte blir en del av den ena skall bli Void. "<Z-Gryphon> som är en slags stor skala, apokalyptisk version av "I            är vad jag äter. ":)
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Liiwi> udp - universal släppa av en duva
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Lilo> Jag har alltid velat ha en webbplats med en stor bild av en morot på det
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Bdale> Bdale är en sammandragning av Barksdale.<Lo-lan-do> Hm. Det är definitivt inte något jag någonsin kommer ihåg.<Lo-lan-do> besvärad om jag kallar dig Wensleydale istället?
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Luca> och de som säger: fiberkablar har en minsta böjningsradie och       pull spänning? bah! *ryck*<CULus> DET ÄR FIBER DU FREAKS: P<Luca> cULus, du Hoser, det är fiber. jag blir tvungen att komma över       berg och ge dig en wedgie?
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Maswan> Joy: Låter gaffel katt! :)<Maswan> Joy: föreställa sig en stor högaffel och en död kattunge ovanpå         det .. med blod rann ..
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Mjg59> Damnit. Jag har en månad att skriva en uppsats. detta innebär        faktiskt skriva bitar av kod jag ska tala        handla om.<Asuffield> hitta ett gäng studenter och ge det till dem som en övning<Mjg59> asuffield: Jag är omgiven av ett gäng studenter. Förra gången jag        låt dem röra kod, kom jag tillbaka och fann de hade skrivas        all C ++ koden i C och alla C-kod i C ++<Asuffield> Mwahaha<Mjg59> och bröt Build
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Moshez> vad jag vill om Manoj är hans önskan om enkla och små         lösningar. liknande EMACS. eller DVT.<Manoj> väl, var DVT _supposed_ att vara enkel<Manoj> det bara tog 2 veckor att skriva<Moshez> Manoj: Det krävs en * schema * att förklara vad varje del gör.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Moshez> ok, kommer jag inte gifta Jo-Con-El ko.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> penis skämt är okej i blandat sällskap. VMS är inte !!!
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> ltd: Fine, gå genom livet bara peka och grymta på            vad menar du. Fungerar för Mac-användare.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
revidering 1.17.2.7datum: 2001/05/31 21:32:44; Författare: Branden; tillstånd: Exp; linjer: +1 -1ARRRRGH !! FICK G ** D *** känslan av ett F ******* TEST baklänges!
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend_> Overfiend första lag Förpackningens Kvalitet: Om             ansvarige gillar att stava en del av eller hela sitt namn i             CAPS, kommer paketet att suga.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend_> Intel. Ger dig det banbrytande teknik från 1979             i 22 år nu.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> nyckeln till korrekt uttal franska är att dra            mungiporna ner så långt som de kan möjligen gå,            och sedan stöna som du förstoppad<Overfiend> du verkligen spika vokalljud på det sättet
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<- Overfiend har slutat ( "våga ut för att förstöra märkliga nya                         världar, och äta liv och nya civilisationer ")
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> typ av landskapet som skrattar åt "AWD" fordon och            skickar dem tumlande i raviner
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> Joy: Hej, jag är en skitstövel. Assholes avger motbjudande gas.            Det är vad vi gör.
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> som aj skulle säga, väntar alltid fungerar<Overfiend> antingen vad du vill händer, eller om du dör och kan inte vara            perturbed anymore<Overfiend> problem med denna filosofi är att aj uppriktigt            anser att det
		-- Shawn McMahon on debian-curiosa@l.d.o

%
* Doogie förvandlas till manoj<Overfiend> doogie: småningom, vi alla förvandlas till Manoj<Overfiend> Manoj är Debians järn<Overfiend> slutligen, vi alla förfall till Manoj
		-- Shawn McMahon on debian-curiosa@l.d.o

%
<Overfiend> men titta på franska. Du kan stava varje ord i            deras språk fonetiskt med endast ca 6 bokstäver<Overfiend> 4 konsonanter och 2 vokaler<Overfiend> c, f, r, l. Och vokaler? Tja, är en ljudet du            gör när du har förstoppning, den andra när du har            diarre<Overfiend> vad förväntar ni er från att kosten sniglar och grodor?
		-- Shawn McMahon on debian-curiosa@l.d.o

%
X-Manoj-Positions Advisory: Observera att Manoj Srivastava sannolikt tvivlar    fakta belägen och motsätter sig alla slutsatser i detta meddelande.
		-- Seen in the headers of a mail from Branden Robinson

%
<Sangr> hem är där den högsta bandbredden är
		-- Seen in the headers of a mail from Branden Robinson

%
<Sangr> inga fler perl ... det är deprimerande ...<Sangr> Jag tror perl och jag behöver lite tid från varandra<Sangr> vi gjorde vacker musik tillsammans ungefär ett år sedan ...<Sangr> men tiderna har förändring, bytte vi ..
		-- Seen in the headers of a mail from Branden Robinson

%
<StevenK> Jag kan oftast dämpar de känslor som säger åt mig att krascha          tackla en flicka in i buskarna
		-- Seen in the headers of a mail from Branden Robinson

%
<Wiggy> bwah, vodka i min mus
		-- Seen in the headers of a mail from Branden Robinson

%
<Wiggy> i en fantastisk ny drag jag faktiskt testat upload
		-- Seen in the headers of a mail from Branden Robinson

%
<WiggyWork> 3990 N 15 april söta flickvän (45) Erotiska Amateur Girlfriends<WiggyWork> Jag var inte medveten om att du hade professionella flickvänner samt
		-- Seen in the headers of a mail from Branden Robinson

%
Dock är min entusiasm för det modulära träd mildras av vissa delar avdet inte existerande.framtid X
		-- Daniel Stone on debian-{x,devel}, commenting on the

%
Har hon tror att vi vill bara sitta målning debian virvlar runt på vårtånaglar?
		-- Erinn Clark, referring to the Debian-women project

%
modconf (0.2.37) stabil instabilt; brådskande = medium  [...]  * Eduard Bloch:    - Fast Make brutit Marcin Owsiany ett tag sedan. Standardmanual      har skrivits över med polsk översättning. Jag undrar fortfarande varför      ingen lade märke till detta innan. Stänger: # 117.474  [...]
		-- Eduard Bloch <blade@debian.org>  Sun, 28 Oct 2001 12:53:27 +0100

%
<| Ryan |> Jag använder inte deb<Netgod> u fattige<Koppla> netgod: heh<Kingsqueak> apt-get install uppgifts p0rn
		-- Eduard Bloch <blade@debian.org>  Sun, 28 Oct 2001 12:53:27 +0100

%
(Det är en gammal Debian tradition att lämna åtminstone två gånger per år ...)
		-- Sven Rudolph

%
<Joey> Gorgo: * lol *<Gorgo> joey: Vad är så roligt? :)<CULus> shh, känguruunge förlorar all sanity från brist på sömn<CULus> ja joey, mycket roligt "<CULus> Humor honom:>
		-- Seen on #Debian

%
* SynrG konstaterar att antalet konfigurations frågor att besvara i sendmail  är icke-triviala
		-- Seen on #Debian

%
* JHM undrar vad Joey gjorde att tjäna "Jag skulle bara vilja säga, för att undvika missförstånd,  att Joey regler. "
		-- Seen on #Debian

%
Har människor som kontrollerar Debians webbplats var 5 minuter för att kontrollera det inteförvandlats till en annan? Inte för att jag är en att prata, men vissa människor på allvarbehöver för att få ett liv.
		-- james on #Debian

%
* james skulle vara mer imponerad om netgod magiska krafter kunde stoppa  delar i första hand ...* Netgod konstaterar Debianutvecklare är notoriskt svårt att imponera
		-- Seen on #Debian

%
   * I väntan på 2.10.02 versionen uppdaterats för att patchlevel     +ircu2.10.01+.config6-7.config7-8.lgline3.iwho.limit.glibc.motdcache2.trace.whois1-2.config8-9.statsw.sprintf2-3.msgtree2.memleak1-2+.msgtree2-3.gline8-9.gline9-10.invite2.rbr.stats.numclients.whisper.whisper1-2.stats1-2.nokick1-2.chroot.config9-11.snomask7-8.limi+t1-3.userip1-3.userip3-4.config11-12.config12-13.umode2-3.akillsbt.who4-5.kn.kn1-2.freebsdcore2.msgtree3-5.y2k.glibc1-2.rmfunc.msgf+lags2.who5-6.nickchange2.glibc2-3.modeless3
		-- From the annoucement of ircd 2.10.01-3 for Debian GNU/Linux

%
* Joey bör inte skriva ändringsposter i 05:30<Joey> * DFSC gratis cgi bibliotek<Joey> Vad är det? DFSC?<jim> Debians fri programvara mroooooCows
		-- Seen on #Debian

%
<James> missbruka mig. Jag är så lame jag skickade en felrapport till debian-devel-changes
		-- Seen on #Debian

%
<Mörk> äter Depends: cook | äta ute.       Men äter ut är non-free så det är ute.       Och kocken rekommenderar: ren-pannor.
		-- Seen on #Debian

%
Du kommer inte censurera mig genom bugg terrorism.
		-- James Troup

%
<Doogie> Thinking är farlig. Det leder till idéer.
		-- Seen on #Debian

%
<James> Ska vi göra en emacs av ​​apt?        APT - Debian i ett program. Det gör även din tvätt
		-- Seen on #Debian

%
Debian är som Suse med yast avstängd, bara bättre. :)
		-- Goswin Brederlow

%
Charles Briscoe-Smith <cpbs@debian.org>:  När allt kommer omkring är gzip paket som kallas 'gzip ", inte` libz-bin "...James Troup <troup@debian.org>:  Eh, antagligen eftersom gzip binära inte kommer från  obefintlig libz paket eller existerande zlib paketet.
		-- debian-bugs-dist

%
<Jim> Lemme göra säker på att jag inte slösa tid här ... bcwhite tar bort      pkgs som havent fastställts som har utestående fel svårighetsgrad      "viktig". Sant eller falskt?<JHM> jim: "viktig" eller högre. Sann.<Jim> Då vi är på väg att förlora ftp.debian.org och dpkg :)* Netgod missar dpkg - det var ibland bra<Joey> Vi har fortfarande rpm ....
		-- Seen on #Debian

%
Att överbelastad är ett tecken på en sann Debianansvarige.
		-- JHM on #Debian

%
Det förvånar mig att ingen bygger en kommersiell distribution på Debianännu - är det överlägset mest solida UNIX-liknande operativsystem jag någonsin installerat,och jag har spelat med HP / UX, Solaris, FreeBSD, BSDi och SCO (intenämna OS / 2, Novell, Win95 / NT)
		-- Nathan E. Norman

%
> <Magisk tre suck av överdrift böjning>Den Branden skuggar din magiska suck. Den Branden attackerar dig med enmassa ord! Den Branden missar!
		-- Henning Makholm in <yahsmr7dk9k.fsf@pc-043.diku.dk>

%
Jag tror inte att "Det är bättre än att kasta sig in i en köttkvarn"är en bra motivering för att göra något.<20030905221055.GA22354@doc.ic.ac.uk> på debian-devel
		-- Andrew Suffield in

%
<Overfiend> whew.<Overfiend> Jag behöver verkligen att få lite sömn.<Overfiend> men det var säkert kul att prata gitarrer, politik och lesbiska.
		-- Andrew Suffield in

%
Den som frågade om debian organisation var död inte läsadebian-devel. 66 meddelanden i en dag, och det är inte över. Jag tycker att det ärsvårt att hänga med.
		-- Bruce Perens

%
<Asuffield> fiber i USA är ett sådant skämt. i de civiliserade delarna av             världen, startar DSL * * vid hastigheter där amerikanska fiber låter off<Joshk> asuffield: Australien är en nation full av vildar?<Asuffield> joshk: de har ungefär en 9600 modem mellan hela             jävla land
		-- in #debian-devel

%
<Nobse> bleh ... kväll hade jag en dröm ... någon NMU'ed vim ...         mardröm
		-- in #debian-devel

%
