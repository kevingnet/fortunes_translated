* SynrG konstaterar att antalet konfigurations frågor att besvara i  send är icke-triviala
		-- David Leimbach

%
* james skulle vara mer imponerad om netgod magiska krafter kunde stoppa  delar i första hand ...* Netgod konstaterar Debianutvecklare är notoriskt svårt att imponera
		-- David Leimbach

%
<Sel> behöver hjälp: min första paketet till min leverantör försvinner :-(<Netgod> sel: inte skicka den första, börja med # 2
		-- David Leimbach

%
<James> missbruka mig. Jag är så lame jag skickade en felrapport till        debian-devel-changes
		-- David Leimbach

%
Jag trodde aldrig att jag skulle se dagen där Netscape är fri programvara ochX11 är patentskyddad. Vi lever i intressanta tider.
		-- Matt Kimball <mkimball@xmission.com>

%
<Jim> Lemme göra säker på att jag inte slösa tid här ... bcwhite tar bort      pkgs som havent fastställts som har utestående fel svårighetsgrad      "viktig". Sant eller falskt?<JHM> jim: "viktig" eller högre. Sann.<Jim> Då vi är på väg att förlora ftp.debian.org och dpkg :)* Netgod missar dpkg - det var ibland bra<Joey> Vi har fortfarande rpm ....
		-- Matt Kimball <mkimball@xmission.com>

%
<JHM> överbelastas är ett tecken på en sann Debianansvarige.
		-- Matt Kimball <mkimball@xmission.com>

%
<Overfiend> partycle: jag på allvar behöver en semester från detta paket.            Jag hade faktiskt en dröm om att införa en dum ny bugg            i xbase-preinst går kväll. Det är ett dåligt tecken.
		-- Matt Kimball <mkimball@xmission.com>

%
Skriva icke-fri programvara är inte ett etiskt legitim verksamhet, så ommänniskor som gör detta stöter på problem, det är bra! Alla företag baseradepå icke-fri programvara borde misslyckas, och ju förr desto bättre.
		-- Richard Stallman

%
Microsoft DNS-tjänsten avslutas onormalt när det tar emot ett svartill en DNS-fråga som aldrig gjordes. Fix Information: Kör din DNStjänst på en annan plattform.
		-- BugTraq

%
* Dpkg händer STU ett stort glas vbeer* Joey tar öl från stu, du är för ung;)* Cylord tar öl från Joey, du är för full.* Cylord ger ölet till muggles.
		-- BugTraq

%
Vi folket av Debian GNU / Linux-distribution, för att bilda enmer perfekt operativsystem, fastställa kvalitet, försäkra marknadenmångfald, sörja för gemensamma behov av datoranvändare, främjasäkerhet och integritet, störta monopolist krafter i datornmjukvaruindustrin, och säkrar välsignelserna av frihet till oss själva ochvåra efterkommande, förordnar och upprättar denna konstitution för DebianGNU / Linux-system.
		-- BugTraq

%
"Detta är den element_data struktur för element vars * ELEMENT_TYPE =FORM_TYPE_SELECT_ONE, FORM_TYPE_SELECT_MULT. * / / * * Häckar djupareoch djupare, hårdare och hårdare, gå, gå, oj, oj, Ohhhhh !! * Tyvärr fickryckas där. * / Struct lo_FormElementOptionData_struct. "
		-- Mozilla source code

%
Medan år 2000 (y2k) problem är inte en fråga för oss, alla Linuximplementeringar kommer påverkas av år 2038 (y2.038k) fråga. DeDebian-projektet har åtagit sig att arbeta med industrin i denna frågaoch vi kommer att få våra fullständiga planer och strategi publiceras under första kvartaletav 2020.
		-- Mozilla source code

%
... Där var Stac Electronics när Microsoft uppfann Doublespace? Varvar Xerox och Apple när Microsoft uppfann GUI? Där var ApplesQuickTime när Microsoft uppfann Video för Windows? Där var SpyglassInc. Mosaic när Microsoft uppfann Internet Explorer? Där var Sunnär Microsoft uppfann Java?
		-- Mozilla source code

%
Jag är ledsen om följande låter stridslysten och alltför personliga,men det är min allmänna stil. - Ian Jackson
		-- Mozilla source code

%
"Mitt största problem med RH (och särskilt RH contrib paket) är attDe har inte något liknande vår politik. Det är en av de främsta anledningarnavarför deras paket är så skit och trasig. Debian har lagarbetesidan av att bygga en distributions ned till en konst. "
		-- Mozilla source code

%
"Slackware användare spelar ingen roll. Enligt min erfarenhet, Slackware användareantingen clueless nybörjare som kommer att ha problem även med tjära, eller så är derabiat gör-det-självare som inte skulle installera någon annans förkompileradebinär även om de betalt för att göra det. "
		-- Mozilla source code

%
<XinkeT> "Herre ge mig sinnesro att acceptera det jag inte kan         ändra, mod att förändra det jag kan, och visdom         att dölja kropparna hos de människor jag var tvungen att döda, eftersom de         gjorde mig arg."
		-- Mozilla source code

%
* Dark har förändrat ämne kanalen #debian till: Senare i kväll: Efter  månader av noggrann kylning, är Debian 2.0 tillräckligt slutligen coolt att  släppa lös.
		-- Mozilla source code

%
Jag satt skrattar snidely i min bärbara dator tills de visade mig en dator medLinux. Och oh! Det var som om himlen öppnade och Gud avkunnats enklientsidan OS så vacker, så graciös och så elegant att en miljonMicrosoft utvecklare kunde inte ha uppfunnit det, även om de hade ett hundratalår och tusen lådor med Jolt Cola.
		-- LAN Times

%
Jag satt skrattar snidely i min bärbara dator tills de visade mig en dator medLinux .... Och gjorde denna dator choke? Har det stamma? Gjorde det, ens en gång,säger att detta program har utfört en förbjuden åtgärd och måste stängasner? Nej Och detta är bara på klienten.
		-- LAN Times

%
"Jag tror att de flesta Debianutvecklare är ganska" viljestark "människormed en hög grad av förståelse och en hög nivå av passion för vadde uppfattar som viktigt i utvecklingen av debian system. "
		-- Bill Leach

%
"Egentligen den enda Linuxdistribution jag någonsin använt som passeraderootshell testet ur lådan (hit rootshell vid den tidpunkt då dist ärfrigörs och se om du kan bryta OS med skript därifrån) ärDebian. "
		-- seen on the Linux security-audit mailing list

%
* CULus fruktar perl - språket med valfria fel
		-- seen on the Linux security-audit mailing list

%
<Stu> bör du vara rädd för att använda KDE eftersom RMS kan komma till      Huset och klyva bildskärmen med en yxa eller något :)
		-- seen on the Linux security-audit mailing list

%
"Och jag faktiskt som Debian 2.0 som mycket jag helt moderniserasStand.inst av Linux-system vårt företag säljer och installeras allaav Linux-system på kontoret och här hemma .. "
		-- seen on the Linux security-audit mailing list

%
<Davide> hur skjutningen en politik polispolitik med en politik för att ändra         polispolispolicy
		-- seen on the Linux security-audit mailing list

%
<Mörk> "Låt oss bilda Linux Standard Linux standardisering Association        Styrelse. Syftet med detta forum är att standardisera Linux        Standardiseringsorganisationer. "
		-- seen on the Linux security-audit mailing list

%
<Overfiend> inte kommer att gråta för mig om dina "30 minuters sammanställer" !! jag            måste bygga X uppförsbacke båda hållen! I snön! med bar            fot! Och vi har inte kompilatorer! Vi var tvungna att översätta            C-kod för att Mnemonics själva!<Overfiend> Och jag var 18 innan vi ens hade montörer!
		-- seen on the Linux security-audit mailing list

%
NEW YORK (CNN) - Internetanvändare som tillbringar även ett par timmar i veckan på nätethemma upplever högre nivåer av depression och ensamhet än omde hade använt datornätverk mindre ofta, The New York Timesrapporterade söndag. Resultatet ... överraskade både forskare ochsponsorer, som ingår Intel Corp., Hewlett Packard, AT & T Forsknings- ochApple Computer.
		-- seen on the Linux security-audit mailing list

%
"Vad som är slående är emellertid den allmänna layouten och integrering avsystem. Debian är en verkligt elegant Linux-distribution; Stor omsorg hartagits i utarbetandet av förpackningar och deras placering inomsystem. Det stora antalet paket som finns tillgängliga är också imponerande .... "
		-- seen on the Linux security-audit mailing list

%
Debian Linux är en solid, omfattande produkt och en verklig glädje attanvändning. Det är också bra att engagera sig med Debian kollektiv,vars vänlighet och anda påminner de första dagarna av Internet ochsin känsla av öppenhet och globalt samarbete.
		-- seen on the Linux security-audit mailing list

%
<Flood> kan jag skriva ett Unix-liknande kärnan i perl?
		-- seen on the Linux security-audit mailing list

%
<Flood> netgod: Jag har också en "Evil Inside" T-shirt (w / Intel-logotypen) .. på        baksidan anges: "När uppryckandet kommer, kommer du att ha root?"
		-- seen on the Linux security-audit mailing list

%
<Zarkov> "NT 5.0. Alla buggar och tio gånger kodstorlek!"
		-- seen on the Linux security-audit mailing list

%
<CULus> finns det 150 meg i / tmp dir! KÄRA HERRE
		-- seen on the Linux security-audit mailing list

%
<Toor> netgod: vad har du i din kärna ??? Den kompilerade källa för       drivning av en rymdfärja ???<Spoo> tid att göra en zip driva diskettenheten sedan. om kärnan       spelar passa på att kärnan är en AI
		-- seen on the Linux security-audit mailing list

%
Nu kan jag äntligen förklara för alla varför jag gör detta. Jag fick bara $ 7 värdav gratis saker för att arbeta på Debian!
		-- seen on the Linux security-audit mailing list

%
<Ultima> netgod: Min miniräknare har flera register än x86, och
		-- thats- sad

%
* Boren kastar Matlab över rummet och hoppas att det bryter sig in i ett antal  aproaching oändliga peices
		-- thats- sad

%
"... Det var en mycket snabbare än jag trodde det skulle vara mycket snabbareän NT. Om ytterligare hastighetsökningar görs till servern för den slutligarelease, är Oracle kommer att kunna torka sin åsna med SQL Server ochlämna det tillbaka till M $ medan Oracle administratörer ... migrera sina databaseröver till Linux! "
		-- thats- sad

%
Världsdominans, naturligtvis. Och lättklädda kvinnor. Vem bryr sig omdess tjugo nedan? - Linus Torvalds
		-- thats- sad

%
<Flav> Win 98 Psychic upplagan: Vi ska berätta vart du ska i morgon
		-- thats- sad

%
<Zpx> det är fantastiskt hur "icke-bruten" debian jämförs med slak och rh
		-- thats- sad

%
<Mörk> "Hej, jag är från detta projekt som kallas Debian ... har du hört talas om det?       Ditt namn verkar vara på ett gäng våra grejer. "
		-- thats- sad

%
"I händelse av en percieved brist av projektet ledar #debian ärbefogenhet att vidta drastiska och descisive åtgärder för att korrigera den felaktiga,bland annat genom att inte begränsad till utvisa tjänstemän, apointing nya tjänstemänoch i allmänhet missbruka makt "
		-- proposed amendment to Debian Constitution

%
<Overfiend> vi kallar 2,2 _POTATO_ ??
		-- proposed amendment to Debian Constitution

%
<SirDibos> gör Johnie Ingram hänga här på IRC?
		-- proposed amendment to Debian Constitution

%
* Twilight1 måste hänga sin Mozilla mössa dinosaurie i effigy om  Netscape säljer ut till många förlorare ..
		-- proposed amendment to Debian Constitution

%
<Lux> om MacOS är för datorn analfabeter, då windoze är för      dator masochister
		-- proposed amendment to Debian Constitution

%
<Mörk> cULus: Att bygga en fem meter hög kopia av Empire State       Byggnad med gem är imponerande. Att göra det med förbundna ögon är       eleet.
		-- proposed amendment to Debian Constitution

%
Jag kan bara se det nu: nominering terrorism ;-)        - Manojhaha! Jag nominera Manoj.
		-- seeS

%
<JHM> På något sätt jag har mer respekt för 14 år gamla Debianutvecklare än     14 år gammal certifierad Microsoft Livegen.
		-- seeS

%
<CULus> Ben: Har du solumly svär att läsa upp debian e en gång om dagen och        tillåter inte folk att tro att du är MIA?<Ben> cULus: jag gör så svär
		-- seeS

%
"Jag undrar om detta är den första konstitutionen i mänsklighetens historiadär man måste beräkna en kvadratroten för att bestämma om en rörelsepasserar. :-) "
		-- Seen on Slashdot

%
Detta är lösningen på Debians problem .. och eftersom det enda riktiga sättetatt skapa fler släktingar av utvecklare är att ha barn, behöver vi mersex! Det är en långsiktig investering ... det är själva arbetet som ärtillfredsställande!
		-- Craig Brozefsky

%
<Marcus> dunham: Du vet hur verkliga siffrorna är tillverkade av rationell         tal av ekvivalensklasser av konvergerande sekvenser?<Dunham> marcus: ja.
		-- Craig Brozefsky

%
<CULus> "Hallå?" "Hej baybee" "Är du Johnie Ingram?" "För att jag ska vara        någon "" Ermm .. Säljer ni slink CD? "" Jag älskar slinkies "
		-- Craig Brozefsky

%
<Overfiend> xhost + localhost endast bör göras av personer som skulle            måla deras värdnamn och rot lösenord på en väg, interstate            viadukt.
		-- Craig Brozefsky

%
<JHM> AIX - Unix från universum där Spock har skägg.
		-- Craig Brozefsky

%
<Knghtbrd> Studier visar att forskningen orsakar cancer i 43% av laboratorie           råttor<CQ> knghtbrd- ja, men 78% av denna statistik är avstängda med 52% ...
		-- Craig Brozefsky

%
<STU> apt: buggar<Apt> buggar är dum<Dpkg> apt: är dumma? vad är det?<Apt> dpkg: Jag vet inte<Dpkg> apt: Skönhet är i ögat av öl hållaren ...<Apt> jag redan hade det på det sättet, dpkg.
		-- Craig Brozefsky

%
<Muggles> jag försöker övertyga några Netcoms administratörer jag vet att konvertera          Debian från RH, netgod, men de är DAMN envis<Muggles> varför RH användare så förbannat hårt väg?<Espy> det är hatten
		-- Craig Brozefsky

%
<Doogie> Debian - All kraft, utan den fåniga hatt.
		-- Craig Brozefsky

%
Hur många månader kommer vi att ligga bakom dem [Redhat] med en glibcsläppa lös?"
		-- Jim Pick, 8 months before Debian 2.0 is finally released

%
Syftet med att ha mailinglistor snarare än med diskussionsgrupper är attplacera ett hinder för inträde som skyddar listorna och deras användare fråninvasion av de allmänna outbildade horder.
		-- Ian Jackson

%
De flesta av oss känner att marknadsföring typer som ett farligt vapen - hålla'Em lossas och inlåst i ett skåp, och bara ta ut dem närdu behöver dem för att göra ett jobb.
		-- Craig Sanders

%
<Benc> Cerb: vi prenumererar du att debian-kamp som moderator<Benc> Cerb: listregler är, 1) ingen trevlig e-post, 2) inga ursäkter
		-- Craig Sanders

%
<Teknix> vår lokala telco har erkänt att någon "backas in i en         knappen på en switch "och tog hela ATM-nätet ner<Netgod> förhoppningsvis nu routrar är utformade bättre, så att "nätverket         off "swtich är på baksidan
		-- Craig Sanders

%
<Overfiend> Thunder-: när du får {MessagesLikeThisFromYourHardDrive}<Overfiend> Thunder-: Antingen sätt {TheDriverIsScrewy}<Overfiend> eller<Overfiend> {YourDriveIsFlakingOut BackUpYourDataBeforeIt'sTooLate            Be till Gud }
		-- Craig Sanders

%
<Apt> har det sagts att RedHat är saken Marc Ewing bär på      hans huvud.
		-- Craig Sanders

%
<MrCurious> i kraft av Greyskull<MrCurious> någon berätta för mig förbudet att placera<Sopwith> mrcurious: * .debian.org, * .novare.net<PhilX> * .debian.org. det är jättebra.
		-- Seen on LinuxNet #linux

%
"Vad gör detta berätta? Att om Microsoft var den sista programvaraFöretaget kvar i världen, 13% av den amerikanska befolkningen skulle skurloppisar och goodwill för gamla TRS-80, CPM maskiner och Apple] [ 's innande skulle köpa Microsoft. Det är inte precis en ringande påskrift. "
		-- Seen on Slashdot

%
"Bruce McKinney, författare av Hardcore Visual Basic, har meddelat atthan trött på VB och kommer inte att skriva en 3: e upplagan av hans bok. Debästa citat är i slutet: "Jag behöver inte ett språk som designats av fokusgrupp'."
		-- Seen on Slashdot

%
<Cylord> Skulle det vara acceptabelt att Debians policy om vi satt i ett crontab         som standard in i potatis som mailade bill.gates@microsoft.com         varje morgon med ett e-postmeddelande som läst, "Oroa dig inte, är Linux en         fluga..."
		-- Seen on Slashdot

%
* Overfiend rar som gör en NMU av asclock, där han ändrar helt enkelt  den förlängda beskrivningen till "Om du böja sig och sätta huvudet mellan  benen, kan du läsa ledigt din assclock. "<Doogie> Overfiend: gå till sängs.
		-- Seen on Slashdot

%
<Reed> Det är viktigt att notera att den främsta orsaken det romerska riket       misslyckas är att de inte hade någon begreppet noll ... vilket de kunde inte       testa framgång eller misslyckande i sina C-program.
		-- Seen on Slashdot

%
Sen när har till syfte att debian varit att blidka intressenmassa outbildade konsumenterna? - Steve Shorter
		-- Seen on Slashdot

%
<Joeyh> netgod: er, är dessa 2.2.0 paket 2.0.0pre9 eller har du en        direkt linje med gudarna?<Netgod> joeyh: Jag har den direkta linjen
		-- Seen on Slashdot

%
<_Anarchy_> Argh .. vem dela ut papperspåsar 8)
		-- Seen on Slashdot

%
<Besvärliga> någon runt?<Flav> nej, vi är alla oregelbundna polygoner
		-- Seen on Slashdot

%
<CULus> OH MY GOD INTE en slumpmässig Quote Generator<Netgod> säkert du tänkte det var statisk? hur lama skulle det vara? :-)
		-- Seen on Slashdot

%
Mere icke-existens är en svag ursäkt för att förklara en sak unseeable. Du* Kan * se drakar. Du behöver bara titta i rätt riktning.
		-- John Hasler

%
<Chalky> gcc är den bästa kompressorn någonsin portas till Linux. den kan vridas         12MB av kärnans källkod (och som .debbed) i en 500k kärna
		-- John Hasler

%
<Manoj> I * som * hönan
		-- John Hasler

%
 [] Dogbert [2] Richard Stallman [3] Buffy Summers [1] Manoj Srivastava [4] Inget av ovanstående
		-- Debian Project Leader 1999 ballot

%
<Oryn> någon som vet om det finns en version av dpkg för RedHat?
		-- Debian Project Leader 1999 ballot

%
acme-kanon (3,1415) instabilt; brådskande = låg  * Extra säkerhet för att förhindra operatören lemlästning, stängs: bug # 98765,    bug # 98713, # 98.714.  * Lade manual. stänger: # 98.725.
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
! Netgod: *! Tiden går fort när youre använder Linux! Doogie: *! yeah, oändliga loopar i 5 sekunder.! Teknix: *! Har någon testas på nytt att med 2.2.x?! Netgod: *! ja, 4 sekunder nu
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
* Mörk hälsar LIW med en liten gul groda.* LIW kysser grodan och klockor det omvandla en vacker nörd  flicka, tar henne ut till glass, och lever lyckligt för evigt efter  med henne<Mörk> LIW: Umm det är för sent att få grodan tillbaka?
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
* CULus anser att vi bör gå till mässor och se hur många människor vi  kan döda genom att kasta Debian-cd på dem
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
<Mörk> "Ja, din ära, har jag RSA krypteringskoden tattood på min        penis. Skall jag visa juryn? "
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
<Knghtbrd> ni är alla vansinniga.<Joey> riddare: säker, det är därför vi arbetar på Debian.<JHM> Knghtbrd: komma i kontakt med din inre galning.
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
<CULus> Saens visar inte mindre än 3 TCP / IP-buggar i 2.2.3
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
<Mercury> alexsh: Var / MYCKET / cairful, kan du, om din otur, steka din          moderkort ..<Knghtbrd> Mercury - låter kul
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
<Rcw> mörk: Caldera?<Knghtbrd> rcw - det är inte en fördelning, det är en förbannelse<Rcw> Knghtbrd: det är en förbannat fördelning
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
Programvaran är som sex, det är bättre när det är gratis. - Linus Torvalds
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
<Mörk> Knghtbrd: Vi har massor av whate.<Knghtbrd> mörk - I Debian? Hell yeah vi gör!
		-- Wile E. Coyote <genius@debian.org>  Sun, 31 Jan 1999 07:49:57 -0600

%
Jag gjorde det bara för att gör dig arg. :-P
		-- Branden Robinson in a message to debian-devel

%
Programvaran krävs Win95 eller bättre, så jag installerade Linux.
		-- Branden Robinson in a message to debian-devel

%
10) Det finns ingen 10, men det lät som ett bra läge :)
		-- Wichert Akkerman

%
Eric Raymond: Jag vill leva i en värld där programmet inte suger.Richard Stallman: All programvara som inte är fri suger.Linus Torvalds: Jag är intresserad av gratis öl.Richard Stallman: Det är okej, så länge jag inte behöver dricka det. jag                   inte gillar öl.
		-- LinuxWorld Expo panel, 4 March 1999

%
Jag är inte en sansade personen ... - Bruce Perens
		-- LinuxWorld Expo panel, 4 March 1999

%
Personligen tror jag inte ofta talar om social bra eftersom när jag hör andrafolk pratar om social bra, det är då jag når min revolver.
		-- Eric Raymond

%
Om vi ​​vill ha något trevligt att få född i nio månader, sedan sex måstehända. Vi vill ha den typ av sex som är acceptabelt och roligt för bådemänniskor, inte den typ där någon få skruvas. Låt oss få några tvärbefruktning, men inte någon få skruvas.
		-- Larry Wall

%
Vi vet alla Linux är stor ... det gör oändliga loopar i 5 sekunder.
		-- Linus Torvalds

%
JA! JA! JA! Oh, ja! (Ooops, jag låter som Meg Ryan ;-)
		-- Ian Nandhra

%
<Knghtbrd> Om jag börjar skriva uppsatser om fri programvara för Slashdot,           vänligen skjuta mig.
		-- Ian Nandhra

%
<RoboHak> hmm, lunch låter som en bra idé<Knghtbrd> skulle smaka som en bra idé också
		-- Ian Nandhra

%
P.S. - Jag är på väg * detta * nära till att köra runt i serverrummet med enpar bultsaxar, och en stor träklubba, skrattar som en galning ochskär allt kan jag passa bultsax runt. och whacking attsom jag inte kan. så om jag verkar halv osammanhängande, eller bara verkligen * verkligen * otäckibland, förlåt mig. stress är ingen vacker sak. }; P
		-- Phillip R. Jaenke

%
Varje företag klagar Microsofts affärsmetoder är helt enkelt enrosenbuske. De ser vackra och luktar trevligt. När en lycklig företag dethronesMicrosoft de kommer att kasta sina kronblad att exponera taggar under. entagg med något annat namn skulle skada så mycket.
		-- Phillip R. Jaenke

%
Något måste görasDetta är någotDärför måste detta göras
		-- The Thatcherite Syllogism

%
<Knghtbrd> xtifr - akta oss för james när han är utanför sin medicin =>
		-- The Thatcherite Syllogism

%
Likgiltighet kommer säkerligen att vara undergång mänskligheten, men vem bryr sig?
		-- The Thatcherite Syllogism

%
Underskatta aldrig kraften i mänsklig dumhet.
		-- Robert A. Heinlein

%
Guld, n .:  En mjuk formbar metall relativt sällsynta i distributionen. Den bryts  djupt i jorden fattiga män som sedan ge den till rika män som omedelbart  begrava tillbaka i jorden i stora fängelser, även om guld inte har gjort  något till dem.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
* Lilo förklarar härmed OPN en virtuell smärta i röven :)
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
"De är både företag - om du har gett dem tillräckligt med pengar, jag ärsäker på att de kommer att göra vad fan du frågar: -> "
		-- David Welton

%
"Du har rätt att inte vara en skitstövel. Om du ger upp denna rättallt du säger och gör här kommer att hållas mot dig. Om du inte kanråd att sluta vara en skitstövel sedan någon kommer att utses att sparkaer härifrån. "
		-- Your rights as an irc addict

%
* Simunye är så glad att hon har sina mödrar genens<Dellaran> du bättre ge tillbaka dem innan hon missar dem!
		-- Your rights as an irc addict

%
<Iambe> lura de intellegent människor på planeten är inte lätt
		-- Your rights as an irc addict

%
Kalifornien, n .:    Från latin "calor", som betyder "heat" (som på engelska "kalori" ellerSpanska "caliente"); och "fornia" "för" samlag "eller"otukt." Därför: Tierra de Kalifornien, "landet av hett sex."
		-- Ed Moran

%
* Caytln slår Lisa<Caytln> catfight: P<LisaHere> Se den flicka, jag gillar det.<LisaHere> :)<Caytln> siffror: D
		-- Ed Moran

%
<MFGolfBal> rit / Ara: Det är något riktigt dement om UNIX            underkläder...
		-- Ed Moran

%
X Window System:  Standarden UNIX grafisk miljö. Med Linux, är det vanligtvis  XFree86 (http://www.xfree86.org). Du kan kalla det X, XFree, X  Window System, XF86, eller en mängd andra saker. Kalla det "XWindows" och  någon kommer att smälla dig och du kommer att ha förtjänat det.
		-- Ed Moran

%
<Knghtbrd> "De samlare valuta är offline." "Jag omdirigering men           de sekundära kopplingar. Om vi ​​omarbeta fas grenrör vi           bör kunna använda plasma spolen matrisen för att manuellt           lansera en ny ostliknande spinoff-serien. "* ShadwDrgn suckar<Fas> du lämna mina grenrör ensam<Fas>!
		-- Ed Moran

%
* Turken tänker små barn är helt bedårande ... especialyy när  de är någon annans.
		-- Ed Moran

%
* Overfiend suckar<Overfiend> Netscape suger.<Overfiend> Det är ett korthus som vilar på en bädd av kvicksand.<Espy> under en jordbävning<Overfiend> i en tornado
		-- Ed Moran

%
<SilverStr> medieetik är en oxymoron, likt Jumbo räkor och            Microsoft Works.<MonkAway> inte tala NT Security
		-- Ed Moran

%
<Silvrbear> Oxymorons? Jag såg en igår - broschyren på "Taco Bell            Näringsinformation "
		-- Ed Moran

%
* Knghtbrd släpper ett par dubbla pipa snurf vapen och täcker  jesus med snurf dart<Jesus> meany: P
		-- Ed Moran

%
<Jgoerzen> doogie: du låter mycket instabil :-)<Knghtbrd> jgoerzen - han är.* Doogie bops Knghtbrd<Knghtbrd> se? Ta till våld = D
		-- Ed Moran

%
Jag har också varit ett stort Unix fan ända sedan jag insåg att SCO var inteUnix. - Dennis Baker
		-- Ed Moran

%
<Dracus> Ctrl + Alt + Kommando + P + R<Knghtbrd> dracus - gudar! Det är värre än EMACS!<LauraDax> hehehehe<Dracus> inte fråga vad som gör: P
		-- Ed Moran

%
<Iambe> du inte är en galning<Knghtbrd> Du uppenbarligen inte känner mig väl nog ännu. =>
		-- Ed Moran

%
* Aj tror Kb ^ Zzz borde plocka olika saker att drömma om än   allmänna resolutioner och politiska förändringar.<Kb ^ Zzz> aj - berätta om det, är detta ett dåligt tecken
		-- Ed Moran

%
<Crow_> hmm, finns det en --now-dammit alternativ för exim?
		-- Ed Moran

%
<DarthVadr> Kira: BLI den mörka sidan, unge.<Kira> darth, jag * är * den mörka sidan.
		-- Ed Moran

%
<Netgod> Fëanor: u har ingen aning om djupet av stupidty av amerikansk lag
		-- Ed Moran

%
Den som sticker ut i mitten av en väg ser ut roadkill för mig.
		-- Linus Torvalds

%
<Lilo> "Vänligen respektera IMMATERIALRÄTT!"<Lilo> "Vänligen visa intellekt." ;)
		-- Linus Torvalds

%
<Knghtbrd> Fëanor - licensfrågor är viktiga. Om vi ​​inte titta på vår           åsnor nu, någon ska komma och bita oss senare ...
		-- Linus Torvalds

%
"Nu ska vi döda dig."
		-- Linus Torvalds

%
* Knghtbrd kan redan föreställa: "Subject: [AVSIKT ATT FÖRBEREDA föreslå   ARKIVERING AV felrapport] stavfel i policydokumentet "
		-- Linus Torvalds

%
<Netgod> heh brinner ett hopplöst fall, som det korrekta uttalet av         "smycke"<Netgod> ge upp :-)<Salvia> och den korrekta stavningen av "färg" :)<Benc> heh<Salvia> och aluminium<Benc> eller kärnvapen<Salvia> du threating mig yankee?<Salvia> bara orsak vi inte har bomben ...<Benc> backa ya gul mage
		-- Linus Torvalds

%
<LauraDax> sett Gud<Tabi-> LauraDax, jag minns inte att se "gud"
		-- Linus Torvalds

%
<Kira> är ett kirurgiskt krig där du går ge de utländska trupperna näsa jobb?
		-- Linus Torvalds

%
<Xtifr> Athena Desktop Environment! I era hjärtan, du * vet * det är        rätt val! :)* Knghtbrd THWAPS xtifr
		-- Linus Torvalds

%
<Knghtbrd> shaleh - orena är bara konstigt.<Espy> heh, är oren sval<Knghtbrd> Espy - och konstigt.<Espy> ja, konstig alltför
		-- Linus Torvalds

%
<Xtifr> direkta hjärnimplantat :)<Knghtbrd> xtifr - yah, sedan använda datorer skulle faktiskt kräva någon           av dessa idioter att tänka!<Knghtbrd>;>
		-- Linus Torvalds

%
<Knghtbrd> Overfiend - BTW tar när vi har upptäckt X hela 1,4 GIGS           att bygga, är du villig erkänna att X är bloatware? =><Overfiend> KB: det finns en 16 halv minut lucka i mitt svar<ACF> knghtbrd: bevis för att X är endast * 2 * värsta fönster      systemet;)
		-- Linus Torvalds

%
<LIW> fan, börjar den autonoma musrörelser vanligtvis efter jag använder en      musknapp<Wichert> inte använder en musknapp då :)<LIW> ja, rätt :)
		-- Linus Torvalds

%
<Knghtbrd> du vet, behöver Linux ett plattformsspel huvudrollen Tux<Knghtbrd> ganska Super Marioish, men med Tux och saker som liten cyber           buggar och borgs och sånt ...<Knghtbrd> Och du måste hoppa förbi billgatus och träffa nyckeln för att släppa honom           i lava och sedan se en kille som ser ut som en RMS           eller någon säga "Tack för att rädda mig Tux, men Linus           Torvalds är i ett annat slott! "
		-- Linus Torvalds

%
<Thoth_> Ja, men det är därför det är numrerade 2.3.1 ... det är för dem av oss         som saknar NT-liknande uptimes
		-- Linus Torvalds

%
<Shinobi> Det finns värre saker än Perl .... ASP kommer att tänka
		-- Linus Torvalds

%
* M2 stirrar på skärmen ... det ser ut som en hamburgare ...<Knghtbrd> m2 - det är ett dåligt tecken
		-- Linus Torvalds

%
<Knghtbrd> Låt den Manoj kalla procmail "ynkliga"
		-- Linus Torvalds

%
<Crow-> Manoj: ja, jag kan inte förstå saker som "s / 3 # $% ^% {]] [@ f245}"<Manoj> Crow: Det är inte riktigt lagligt ;-)<Knghtbrd> Manoj - hur skulle man göra "s / 3 # $% ^% {]] [@ f245}" laglig           i alla fall? (Och vad skulle det göra? Hehe)<Manoj> Knghtbrd: Du måste avsluta s /// uttryck.<Knghtbrd> åh, det är allt?
		-- Linus Torvalds

%
<Kira> Ada, det enda språk skrivs till milspec.<Mikster> <ryser>
		-- Linus Torvalds

%
<Benc> -Includemeny ../../debian/el33t.h<Benc> sendmail bygga ... konstigt rubriknamn :)<Isildur> hahaha* netgod laffs<Netgod> Benc: kan u berätta jag brukade hålla sendmail? : P<Benc> heh :)
		-- Linus Torvalds

%
<Fas> nej ... jag musn't ha mer kaffe !!! ;)<Simunye> säker yu göra Fas :)<Fas> du verkligen vill mig studsar taket?<Simunye> Yesh :)<Kira_> studsar taket är gewd<Fas> ok, det var en dum fråga<Kira_> det splatting på golvet som är problemet.
		-- Linus Torvalds

%
<Kensey> RMS för President ???<RelDrgn> ... eller ESR, vill han ett nytt jobb;)
		-- Linus Torvalds

%
Åh nej, inte igen.
		-- Manoj Srivastava

%
<Knghtbrd> Visst, RMS är en fanatiker, jag förnekar inte detta. Jag ska även säga           Han är en kunglig smärta i röven för det mesta. Men han är           ännu oftare rätt än inte, och han förtjänar en viss nivå av           kredit och respekt för sitt arbete. Vi skulle inte vara här i dag           utan honom.
		-- Manoj Srivastava

%
<Espy> i morgon kommer det att finnas en stor störning i arbetskraften
		-- May 18, 1999

%
Jag är dyslektiker av Borg. Förbered dig på att få din röv laminerade.
		-- May 18, 1999

%
<NeonKttn> Jag hade en vän hålla mig i hennes garderob under highschool beacuse I           skulle inte tro att hennes pojkvän visste om förspel ...<NeonKttn> I shoulda fört popcorn. :)
		-- May 18, 1999

%
<Knghtbrd> hardcopy är för wussies<Topher> dator programförteckningar .... nästa, på Hardcopy
		-- May 18, 1999

%
<Kceee ^> Jag hatar användare<Knghtbrd> du låter som en sysadmin redan!
		-- May 18, 1999

%
<Change_m2> Will LINUX någonsin köra skivat bröd som # 1 prestation            mänskligheten?
		-- May 18, 1999

%
<APH> manoj går muttrar på felrättning korståg! woo woo!<Knghtbrd> manoj gick nötter för länge sedan. men felrättning är cool =>
		-- May 18, 1999

%
<Rcw> dessa till synes-bakterier liknande multi maskar kommer ut ur      Microsofts BackOrifice<Rcw> det är backoffice logo
		-- May 18, 1999

%
* Simunye är på en oc3-> Oc12<Daem0n> simmy: bita mig. :)<Simunye> demonen: okej :)
		-- May 18, 1999

%
<Overfiend> lilo: Nåväl, är du förmodligen en ansvarig tänkare.            Välkommen till en mycket liten klubb.<Lilo> Overfiend: välkomna mig när du går :)
		-- May 18, 1999

%
I grund och botten vill jag att folk ska veta att när de använder binär bara moduler,Det är deras problem. Jag vill att folk ska veta att i deras ben, och jagvill ha det ropade från hustaken. Jag vill att folk ska vakna upp i enkallsvett varje gång på ett tag om de använder binär enbart moduler.
		-- Linus Torvalds

%
* Wichert_ föreställer mästare utan MTA<James> Wichert: EHM? som kan hindra peformance av BTS: p
		-- Linus Torvalds

%
<Gecko> Hmm ... jag undrar vad separerar Debian från resten av        Linux-distributioner.<Knghtbrd> gecko - Vi inte suger<Gecko> Knghtbrd: du behöver inte säga att när man hanterar en massa människor        Från dessa distributioner<Knghtbrd> gecko - punkt.
		-- Linus Torvalds

%
På grund av modellen stängd källkod utveckling XFree det är omöjligtatt stödja eller ens spekulera om, funktioner pre- eller betaversionerav XFree.
		-- Marcus Sundberg

%
>> Jag vet inte riktigt ser bibel-kjv-text som ett tekniskt dokument,>> Men ... :)> Det är en handbok - för att leva.Men det inte har uppdaterats på länge, skulle många säga att det ärtyvärr föråldrad och uppströms ansvarige inte svarar på hanse-post. :-)        - Branden Robinson, Oliver Elphick och Chris Waters i en           meddelande till debian-policy
		-- Marcus Sundberg

%
<Knghtbrd> Jag kan tänka mig massor av människor som behöver user = ID10T någonstans!
		-- Marcus Sundberg

%
<Slashdot> min amerikanska geograpy är usel ... lol<Knghtbrd> så är min och jag bor här
		-- Marcus Sundberg

%
Moonchild utan en åsikt? Satan skridskor till jobbet i morgon!
		-- Brett Manz

%
<Knghtbrd> Jag vill verkligen inte mycket alls ... Bara ett vänligt ord, en           attraktiv kvinna, och Obegränsad bandbredd !!
		-- Brett Manz

%
<Knghtbrd> Om vi ​​är båda rätt (jag gissar vi) Jag är inte glad.* Minupla händer dig drift of the Year.
		-- Brett Manz

%
Förra gången jag hade intim kontakt med en annan människa var snarare ensmärtsam upplevelse ... jag hellre velat det ...;)
		-- Brett Manz

%
<Apple_IIe> någon sett min 80 kolonn kort?
		-- Brett Manz

%
<Slackware> uh oh, vad har jag började :)<Debian> rofl ... distro nick krig.* Slackware väntar bara för / nick Gnome, / nick KDE, och sedan andra världskriget 4   att bryta ut<WinNT>: oP<OpenBSD> <anka><PalmOS> :)<Slackware> no'one skulle våga / nick RedHat<Tru64> mew.
		-- Brett Manz

%
<Crow-> im fcucking druk* Knghtbrd ser att logga allt Crow- säger i kväll ...<MrBump> heheh<MrBump> Han sade att han skulle gifta sig med mig! helvete!!<Crow-> dude inget sätt<Knghtbrd> MrBump - han inte som berusad<MrBump> Knghtbrd: Jag krossade: o)
		-- Brett Manz

%
<Knghtbrd> aggh!<Knghtbrd> GÖR DET ATT STOPPA!<Knghtbrd> GÖR DET ATT STOPPA !!
		-- Brett Manz

%
<Knghtbrd> RoboHak - okej, plåstret inte bruten, men min hjärna           uppenbarligen är<Wc> det är inget nytt (;<Knghtbrd> wc - hysch.<Knghtbrd> =>
		-- Brett Manz

%
<DPG> amerikaner är Yahoo ....<Xtifr> Californians ännu weirder<Knghtbrd> xtifr har en punkt ...
		-- Brett Manz

%
* Woot ler serenely.<Woot> Jag vill inte verka över angelägna om att få in knghtbrd s       siglist.
		-- Brett Manz

%
<CULus> dhd: R du en del av hemligheten debian overstructure?<DHD> nej. det är ingen hemlighet debian overstructure.<Kosmiska partiklar> men nu när någon tog upp det, låt oss börja en            :-)<Knghtbrd> kosmiska partiklar - varför inte, låter som ett roligt sätt att tillbringa           eftermiddag = D
		-- Brett Manz

%
<Xtifr> du behöver inte vara galen för att arbeta här .... oh vänta, ja du gör!        :)
		-- Brett Manz

%
* O-o alltid som debmake eftersom han visste exakt vad det skulle göra ...<Ibid> o-o: ni skulle ;-)
		-- Brett Manz

%
2.3.1 har släppts. Folks ny på detta spel bör komma ihåg att2.3. * Utgåvor är utvecklings kärnor, med inga garantier för att deinte kommer att orsaka systemet att göra hemska saker som korrupta dessdiskar, fatta eld, eller börja köra Mindcraft riktmärken.
		-- Slashdot

%
do {    :} While (HELL_FROZEN_OVER!);
		-- Slashdot

%
0 7 * * * echo "... Linux är bara en modefluga" | post billg@microsoft.com -s = "Och kom ihåg ..."
		-- Slashdot

%
<Hop> kb: Jag kräver integritet och ärlighet hos dem som jag gör affärer med<Hop> jag vet mina krav är orimliga, men en kille kan drömma, kan inte han?
		-- Slashdot

%
<Jgoerzen> stu: ahh den maskinen. Tror du inte att något som heter           Stallman förtjänar att vara en Alpha? :-)<Stu> jgoerzen: nej, faktiskt, jag skulle prolly vara mer benägna att nämna 386      med 4 meg RAM och en 40 meg hårddisk Stallman.<Stu> med en stor fet fall som gör massor av buller och skramlar golvet* Knghtbrd faller till golvet håller sina sidor skrattar<Stu> och ..<Stu> dubbel höjd hårddisk
		-- Slashdot

%
Klingon funktionsanrop inte har "parametrar" - de har argument "
		-- and they ALWAYS WIN THEM.

%
* Knghtktty inte kommer att fråga hur zucchini kom in i diskussionen ...
		-- and they ALWAYS WIN THEM.

%
<Knghtbrd> Ämne: [GR FÖRSLAG] Ska vi rösta om triviala frågor?
		-- and they ALWAYS WIN THEM.

%
<Woot> Sätt * att * i dig .sig och rök det, Knghtbrd.<CULus> Du vet att han kommer att läsa detta:><Woot> heheheheh.
		-- and they ALWAYS WIN THEM.

%
"Som ni resa genom livet ta en minut då och då för att ge entrodde för andra kolleger. Han kan rita något. "
		-- Hagar the Horrible

%
<Knghtbrd> Okej, du folk har börjat prata om BSDM tillämpningar av           nätverkshårdvara ... Jag tror att jag ska springa iväg och göra något nyttigt           och Debianish och hålla sig borta från den här ...<Knghtbrd> (för en förändring)
		-- Hagar the Horrible

%
<Knghtbrd> mariab - tror inte att Debian har inte haft några mycket dum och           uppenbara buggar innan<Knghtbrd> naturligtvis vi brukar fixa vår innan vi släpper = D
		-- Hagar the Horrible

%
<Knghtbrd> mariab - Jag är en Debianutvecklare. Red Hat är "fienden" eller           något som jag antar .. Still, type-casting RH användare som           idioter eller deras fördelning så fullständigt bryts av standard           är fullständig och total FUD.
		-- Hagar the Horrible

%
>> Men IANAL, naturligtvis.>> IANAL heller. Min son är, men om jag frågade honom jag kan få ett svar jag> Vill inte höra."Här är min faktura." ? = D
		-- Hagar the Horrible

%
> Ok, jag ser att du vet vad du gör :-)Antingen det eller jag har blivit ganska bra på att fejka det.
		-- Hagar the Horrible

%
<Wichert> 8:00 är en ungoldly timme att vara vaken :)* Gorgo blir oftast upp vid 11:00
		-- Hagar the Horrible

%
Det finns ingen Cabal.
		-- Hagar the Horrible

%
<_Anarchy_> ACF: kanske April 1 nästa år slashdot behöver köra "Rob Malda            accepterar nya jobb som chef för Debian-projektet "8)
		-- Hagar the Horrible

%
* Netgod öppnar sin postlåda och omedelbart vill han hadnt
		-- Hagar the Horrible

%
<Frogbert> det är svårt att vara en lesbisk withoutn bröst ... folk fattar           du på allvar
		-- Hagar the Horrible

%
Kanske Debian är oroad mer om teknisk kompetens snarare änanvändarvänlighet genom att bryta programvara. I det förstnämnda kan vi excel. isenare måste vi medge fältet till Microsoft. Gissa var jag vill gåi dag?
		-- Manoj Srivastava

%
* PerlGeek är verkligen en utomjording* Knghtktty tror PerlGeek
		-- Manoj Srivastava

%
<Netgod> min klient har ägts allvarligt<Netgod> här killen fick rot, sprang Paketsniffare, installerade .rhosts ochbakdörrar, sätta en helt ny dir i kallas / lib / "", som har enkomplett uppsättning smurfing och döda verktyg<Netgod> den enda misstag var inte att ta bort loggfilerna<Netgod> fråga är hur var rot hackat, och att jag kunde berätta u<Netgod> det är, naturligtvis, inte en debian låda* Netgod noterar debian rutan är den enda kvar orört av hackare
		-- wonder why

%
* joeyh cvs begår sin hemkatalog. aaaaaa<Drow> eeeeeeek<Drow> joeyh: Det är helt enkelt ont. Period.
		-- wonder why

%
<Kethryvis> Gruuk: UFies är utöver den mänskliga rasen :)
		-- wonder why

%
Jag slutade för länge sedan för att försöka hitta något i bugg listan över dpkg.Vi ska köra för en post i Guinness rekordbok.
		-- Stephane Bortzmeyer

%
<Ahzz_> i figured 17G oughta vara tillräckligt.
		-- Stephane Bortzmeyer

%
<N3tg0d> har / usr / bin / emacs satts i / etc / shells ännu? : P
		-- Stephane Bortzmeyer

%
* Joeyh utnyttjar Netscapes fantastisk förmåga att krascha för att stänga        10 fönster med en enda knapptryckning<Joeyh> nu det är framsteg!<Knghtbrd> Bussfel =>
		-- Stephane Bortzmeyer

%
<Ordlekar> Du mäter dina vibratorer i "tecken per sekund"? jag hardåliga nyheter för dig, C90, du har onanerar med enmatrisskrivare.
		-- Stephane Bortzmeyer

%
Hej! Jag är en .signature virus! Kopiera mig i din ~ / .signature att hjälpa mig Sprea =d!
		-- Stephane Bortzmeyer

%
* Knghtktty viskar gulligt nonsens till Thyla (saker om kompilatorer och            grafik och uppgraderingar RAM och stora hårddiskar ...)<Thyla> oooooooooOOOOOOOOOO<Infinitas> Knghtktty: det är positivt pornografiskt ...* Thyla går ut i anfall av extas ...
		-- Stephane Bortzmeyer

%
<Sanaya> ni är alla sjuka! sjuk sjuk sjuk jag säga ya;)
		-- Stephane Bortzmeyer

%
* Bma är en ryck* Knghtbrd är en Knghtbrd* DHD är också ett ryck* Espy är ont* Knghtbrd tror Espy
		-- Stephane Bortzmeyer

%
* Bma undrar om detta kommer att göra Knghtbrd .sig
		-- Stephane Bortzmeyer

%
Techical lösningar är inte en fråga om att rösta. Två lagstiftning i USAstater nästan beslutat att värdet av Pi vara 3,14, exakt. folkomröstninggör inte en korrekt lösning.
		-- Manoj Srivastava

%
<Aj> <Knghtbrd> ökningen i spänning i hela världen (vilket framgår av brott<Aj> och allt) under denna tidsperiod ser ut ungefär som Linux<Aj> tillväxt sedan 1993<Aj> `` Linux kopplade till världs brott epidemi !! ''
		-- Manoj Srivastava

%
<Teller> där är jag och vad jag gör i denna handbasket?
		-- Manoj Srivastava

%
Eftersom denna databas inte används för vinst, och eftersom hela verk är intepublicerat, faller det under fair use, som vi förstår det. Emellertid, om någonhalf-assed idiot beslutar att göra en vinst på detta, måste dedubbelkolla allt ...
		-- Notes included with the default fortunes database

%
Det finns ingen snooze-knappen på en katt som vill ha frukost.
		-- Notes included with the default fortunes database

%
Ämne: Bug # 42432: debian-policy: Förslag till CTV för Utkast till Bevis påKoncept för Förslag Förslag till Förslag till CTV till CTV att besluta omett förslag till CTV för CTV på huruvida vi shoud har en CTV på/ usr / doc till / usr / share / doc övergång nu eller senare.
		-- Ed Lang

%
<Knghtbrd> Det är en styrkula för en<Wichert> så det inte är en gnagare<Wichert> det är en skit med en boll som sticker ut<Wichert> som du smeka ständigt
		-- Ed Lang

%
* HomeySan väntar på Papa John pizza att visa upp<Ravenos> mm. Papa John.<HomeySan> förhoppningsvis de skickar söta leveranschaufför<Ravenos> de inte har det här.<Dr_Stein> varför? Ska du äta föraren istället?
		-- Ed Lang

%
<Netgod> är det mig, eller Knghtbrd snarkning?<Joeyh> de dödade knghtbrd!<Netgod> Kysh: Wichert, gecko, joeyh, och jag är i ett rum som försöker ignorera          Knghtbrd<Kysh> netgod: Knghtbrd är svårt att bortse från.
		-- Ed Lang

%
<Woot> Man vill jag knghtbrd var här för att ta det för hans sig listan.[... Flera timmar senare ...]<Knghtbrd> vet woot mig inte vewy bra, gör han?<Knghtbrd> muahahahaha
		-- Ed Lang

%
* Knghtbrd skinn Wichert med NERF dart* Wichert Anteckningar Det finns inga ICBM nerfs ännu och ignorerar kngtbrd<Knghtbrd> Wichert - bara vänta, efter att ha sett NERF Gatling vapen, ICBMs           är inte långt borta (bara pumpa förbannade sak för en timme eller två           är allt...)
		-- Ed Lang

%
Operativsystem Installerad:  * Debian GNU / Linux 2.1 4 CD Set ($ 20 från www.chguy.net; priset ingår    skatter, sjöfart, och en $ 3 donation till FSF). 2 CD är binärer, 2 CD    kompletta källkoden;  * Windows 98 Second Edition Upgrade version ($ 136 genom Megadepot.com,    Priset inkluderar inte skatter / frakt). Överraskande, ingen källkod    ingår.
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
Stjäla detta slogan. Jag gjorde.
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
<Bfextu> oh noooo fick Knghtbrd är en pistol :)<Doogie> ^^ infoga musik ^^<Knghtbrd> bfextu - o / ~ alla är på flykt o / ~<Bfextu> o / ~ springa iväg, ruuuuun bort från betal-ay-ain o / ~
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
<Mercury> emacs suger, bokstavligen, inte en förolämpning, bara en kommentar att dess          stor nog att ha en märkbar gravitationskraft ...
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
Som en dator, jag tycker din tro på teknik underhållande.
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
* Knghtbrd delar 3 till Chris* variabla undrar vem namnges chris förutom mig<Knghtbrd> variabel - du. =>* Knghtbrd väntar variabel att dramatiskt säga "Jag känner mig så används!"<Variabel> Knghtbrd: :)* Variabel ++<Variabel> :)
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
* Espy funderar en uplad kö som kallas "helvetet" så jag kan göra dupload --to helvetet
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
<Valkyrja> java, hon, ibland vill jag verkligen att smälla dig.<Knghtbrd> Valkyrja - han skulle njuta av det för mycket<Reteo> Valkyrja: yah, gå vidare och göra det ... slå java i cappuccino! :-)
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
<Tali> vara vewwy vewwy qwuiet .. Jag är Huntin wuntime ewwos
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
Red Hat har nyligen släppt en Security Advisory (RHSA-1999: 030-01)omfattar ett buffertspill i vixie cron paketet. Debian harupptäckte felet två år sedan och fast det. Därför versionerbåda, den stabila och den instabila, distributioner av Debian inte ärsårbara för detta problem ..
		-- Bill Stilwell, http://linuxtoday.com/stories/8794.html

%
Först ut - Quake är helt enkelt otroligt. Det låter dig upprepade gånger döda dinchef på kontoret utan att gripas. :)
		-- Signal 11, in a slashdot comment

%
Lucas lag: Bra kommer alltid att vinna, eftersom det onda hyr _stupid_             ingenjörer.
		-- Signal 11, in a slashdot comment

%
* TribFurry bara får skräppost från UCSD ... Jag brukade få e-post från            själv men jag bestämde jag inte gillar mig och slutade prata	    till mig
		-- Signal 11, in a slashdot comment

%
<Rain_work> anteckning på en studentrummet kylskåp ... "till den person som åt innehållet            av behållaren märkt "James" - varning, det var min biologiexperiment "
		-- Signal 11, in a slashdot comment

%
<KatanaJ> Obs på en chem lab kyl "Kylskåpet är inte explosions          bevis".
		-- Signal 11, in a slashdot comment

%
<KnaraKat> DalNet är som Special Olympics i IRC. Det finns en hel del           dreglande goin 'on och alla är en "vinnare".
		-- Signal 11, in a slashdot comment

%
Men modifiera dpkg är omöjligt, och vi har kommit överens om att, bland annat,hålla behoven hos våra användare i spetsen för våra sinnen. Och från enanvändarens perspektiv, något som håller systemet snyggt i det normalafall, och arbetar * nu * är mycket bättre än idealistiska fantasier som enarbets dpkg.
		-- Manoj Srivastava

%
För varje visionen finns en lika stor och motsatt översyn.
		-- Manoj Srivastava

%
<Epsilon3> Knghtbrd, om vi ville ha en lameass anmärkning vi skulle ha sagt:           Hej, neckro
		-- Manoj Srivastava

%
<Tigah _-> Jag har 4gb för / tmp<Knghtbrd> Vad gör man med 4G / tmp? Kompilera X?<Tigah _-> ja
		-- Manoj Srivastava

%
<KnaraKat> Bite mig.* TheOne blir lite salt, fortsätter sedan att knapra på KnaraKat lite         bit....
		-- Manoj Srivastava

%
* Knghtbrd konstaterar han har potatismos för hjärnor kväll<Valkyrie> yum, kan jag ha lite?<Knghtbrd> um ...* Knghtbrd hudar från Valkyrie
		-- Manoj Srivastava

%
<Knghtbrd> joeyh har nu en terminal på soffan?<Knghtbrd> Att killen är fast, svär jag =><Doogie> Knghtbrd: laptop<Doogie> och jag menar inte katterna.
		-- Manoj Srivastava

%
Med tanke på några av de senaste trådarna, de interaktiva diskussioner kanskemåste utföras på duk, i närvaro av en domare, medanbär vadderade handskar. ;-)
		-- Phil Hands

%
<James> men sedan jag använde en Atari, jag var mer sannolikt att vinna på lotteri i        tio länder samtidigt än att få snabbare X
		-- Phil Hands

%
* Joeyh undrar varför alla vill veta hur lång han är<James> joeyh: det hjälper sniper
		-- Phil Hands

%
* Benc undrar varför han har uppgraderats till 3.3.5-1 innan coh X ansvarig
		-- Phil Hands

%
<Delenn> Jag skulle inte göra det genom 24 timmar innan jag skulle skjuta upp         grill och slapping några vänner på barbie.<Spacemoos> Varför skulle du smälla vänner med barbies, brinner kinda kinky
		-- Phil Hands

%
I själva verket .. bygger på denna modell av vad NSA är och är inte ... många avmänniskor som läser detta är medlemmar av NSA ... /. är afterall 'News förNerds ".NSA måndag morgon {vid kaffemaskin):NSA AGENT 1: Hey guys, gjorde du kolla in slashdot under helgen?    AGENT 2: Nej, jag har installerat Mandrake 6.1 och jag coulnd't få darn             PPP-anslutning upp ..    AGENT 1: Tja checka ut ... de är på oss.
		-- Chris Moyer <cdmoyer@starmail.com>

%
Tekniken en constand kamp mellan tillverkare som producerar större ochmer idiotsäkra system och natur som producerar större och bättre idioter.
		-- Slashdot signature

%
knghtbrd: det kan finnas någon sked, men kan du upptäcka sårbarheten ieye_render_shiny_object.c?
		-- rcw

%
<Joy> wow ... enkla matematik visar att Debianutvecklare har stängt mer      än * 31 * * tusen * felrapporter sedan vår BTS existerar!<Joy> som är ungefär 30.999 mer än Microsoft;)
		-- rcw

%
<Knghtbrd> OBS att ovanstående är bara en åsikt och bör inte varaAnses omfatta alla former av fakta. DE           TALARE SÄGER allt och alla. HANTERA DET.
		-- rcw

%
<James> GNOME freaks runt?<Knghtbrd> inte mig, jag är bara ett missfoster
		-- rcw

%
<Madax> ahh<Madax> en samling av nördar ....<Madax> Jag kan luktar det nu
		-- rcw

%
<Knghtbrd> lära sig att älska Window Maker.<Knghtbrd> lite Nextstep är bra för själen.
		-- rcw

%
Varningar: det är GNOME, vara rädd, vara mycket rädd för Depends linje
		-- James Troup

%
<CULus> Hhhmmmmmmmm<cULus> vattensängar för kor<CULus> eleet<Cas> cULus: varför skulle en ko behöver en vattensäng?<CULus> cas: Att vara bekväma varm
		-- James Troup

%
Om du är vad du äter, jag antar att det gör mig en ost danska.
		-- Anonymous

%
<Hop> när du börjar göra bara dumma misstag som är uppenbara, brinner      när du börjar få kompetent<Hop> eftersom du inte göra grundläggande missförstånd misstag<Hop> och brinner * bra * tecken.
		-- Anonymous

%
<Lilo> det är konstigt, när man går på en safari till Afrika för att fånga ett lejon, du       tycker att det är levande och det tar, och sedan döda den<Lilo> när du går på en safari till South Bay för att hitta en Palm Vx, hittar       det döda och ta hem och det tar efter det kommer :)
		-- Anonymous

%
<Lilo> Jag kan läsa den blodiga * manuell * som om det vore något slags       religiösa systemet former av upplysning du kan uppnå beskriva       efter 10 år på ett berg :)
		-- Anonymous

%
Gates lag: Var 18 månader, hastigheten på programvaru halvor.
		-- Anonymous

%
<Knghtbrd> Solver_: lägga till användare som ska jävlas med ljud att gruppera           ljud .. Kontrollera att enheterna är alla grupp ljud (ls -l           / Dev / dsp ger dig den snabbaste indikation om det är sannoliktinställd till höger) och bygga en kärna med ljud stöd för kortet<Knghtbrd> eller eventuellt installera alsa källa och bygga moduler för att           med make-kpkg<Knghtbrd> ELLER (rekommenderas inte) få och installera onda OSS / Linux ont           icke-fria onda binära endast onda förare --- men de är onda.Och nämnde jag att det inte rekommenderas?
		-- Anonymous

%
Jag tror irc kommer inte att fungera om --- vi kör ut ur ämnet utrymme!
		-- Joseph Carter

%
"Pacific Bell kundservice, är detta [..], hur kan jag ge digutmärkt kundservice i dag? ""Hahahahaha !! Det är bra, jag gillar det ..""Um, tack, de gör oss säga det."
		-- knghtbrd and a pacbell rep, name removed to protect her job

%
<Danpat> Omnic: blodiga newzealanders<Omnic> danpat: sätta en strumpa i det<Danpat> heh :)<Knghtbrd> gör narr av .nz'ers är annorlunda --- de är alla konstiga* knghtbrd hudar<Omnic> hrmph
		-- knghtbrd and a pacbell rep, name removed to protect her job

%
<Joy> Flinny: svart crontab magi kinda saker :)<Knghtbrd> Joy: Betyder det människor får dansa naken runt bål           mäss konstiga saker och vifta med sina armar omkring i en dum           sätt?<Rcw> knghtbrd: vad tycker du * tror * människor gör på Novare?
		-- knghtbrd and a pacbell rep, name removed to protect her job

%
<Knghtbrd> * snipsnip *<Rcw> Åh kära, är att ljudet av förmögenhet-databas redigering?<Joy> uh oh<Knghtbrd> Ja =>
		-- knghtbrd and a pacbell rep, name removed to protect her job

%
<Joy> som är en Kludge (TM)<Knghtbrd> Det fungerar (tm)<Joy> AIX fungerar (TM)<Knghtbrd> nej det inte<Knghtbrd> =>
		-- knghtbrd and a pacbell rep, name removed to protect her job

%
"Skillnaden mellan snille och stupidity är att snille har detgränser. "
		-- Albert Einstein

%
<Knghtbrd> Om laddnings någon för brott mot USA: s krypto lagar skulle få           du skrattade utanför domstol, bara "undersöka" dem på orättvist laddning           för förräderi!<Knghtbrd> Tea, någon?<Espy> jag hellre dränka politiker i stället för te :)<Stu> espy: politiker har gälar, duh<ESPY> vesslor inte har gälar
		-- Albert Einstein

%
Om jag har problem med att installera Linux, är något fel. Mycket fel.
		-- Linus Torvalds

%
* Bma_home trevar dig<Bma_home> "oups, fel kanal"<Bma_home> </ acf><Cerb> quit groping mig<Doogie> du vet att du gillar det.<Bma_home> faktiskt, att det var "grope me baby"<Gecko-> röra min son och du dör, bma;)<Doogie> gecko-: men din fru är ok?
		-- Linus Torvalds

%
Läsa handböcker dator utan hårdvaran är så frustrerande som läsningkön manualer utan programvaran.
		-- Arthur C Clarke

%
<Knghtbrd> (tinc)<Espy> (ytitac)<Knghtbrd> (ntinac)<Espy> (det)<Knghtbrd> (i)* Espy konstaterar talar i ACR ^ Winitialisms är skrämmande när den andra sidan  förstår dig
		-- Arthur C Clarke

%
<Knghtbrd> Det är synd äldsta Unix är Y2K kompatibel<| Regn |> synd?<| Regn |> varför, eftersom människor inte kommer att uppgradera förrän 2038?
		-- Arthur C Clarke

%
<Espy_on_crack> "Jag installerade" Linux 6.1 ", inte att göra mig en Unix                guru?"<Benc> Espy_on_crack: nej, måste du installera det två gånger innan du är en       guru ... en gång för att bevisa att du kan göra det, det andra att fastställa saker       din bröt första gången<Espy_on_crack> oh rätt, hur dumt av mig
		-- Arthur C Clarke

%
* Knghtbrd gör ET sak<Knghtbrd> någon fick en tala-n-spell?
		-- Arthur C Clarke

%
<Omnic> annan .sig tillsats
		-- Arthur C Clarke

%
Jag börjar tro att genpoolen kan använda lite klor.
		-- Arthur C Clarke

%
Det är så illa som du tror, ​​och de är ute efter dig.
		-- Arthur C Clarke

%
<Espy> vara försiktig, kan vissa twit citera<Espy> ur sitt sammanhang ...
		-- Arthur C Clarke

%
*** Ämne för #redhat: Redhat är svaret på alla dina problem. Det    kan vara början också!
		-- Arthur C Clarke

%
* Cesarb undrar om mindre än en vecka Carmack kommer att hamna emot i  e-posta en artighet kopia av en version av Quake källa som är fyra  gånger snabbare än vad som gick ut ur hans virtuella händer ...
		-- Arthur C Clarke

%
<Knghtbrd> JHM: Jag sätter inte skalvet i kärnan källa<Knghtbrd> men vi bör sätta skalvet i startdisketterna till en upp           Caldera s Tetris spel ..;>
		-- Arthur C Clarke

%
Vapen dödar inte folk. Det är dessa jävla kulor. Guns bara få dem attriktigt riktigt snabbt.
		-- Jake Johanson

%
<Espy> vi måste dela på i "kärnan" och "wtf användnings-här"
		-- Jake Johanson

%
<Culus-> libc6 är inte nödvändigt: |
		-- Jake Johanson

%
<DHD> finns det en speciell jul pack för skalvet<DHD> där du får vara santa robot på futurama?<Dunham> DHD: det skulle vara en ganska obalanserad spel ...<Knghtbrd> dunham: det är tanken. ;>
		-- Jake Johanson

%
<Knghtbrd> problemet med GNU kodningsstandarder är de antar attalla i världen använder emacs .. Om så vore fallet, gratis           programvara skulle dö eftersom vi alla skulle ha handledsproblemsom RMS av nu och inte längre kunna koda. ;>
		-- Jake Johanson

%
C'mon! politisk protest! sheesh. Var är det anarkistiska anda? ;-)
		-- Decklin Foster

%
Vi har höjt våra normer, så upp din!
		-- Decklin Foster

%
* Woot är nu känd som woot-middag* Knghtbrd strör lite salt på woot<Knghtbrd> Jag har aldrig haft en woot innan ... Hoppas de smakar bra<Woot-middag> noooo!<Woot middagen> äter inte mig!* Knghtbrd bestämmer han inte vill ha en middag som talar till honom ... hehe
		-- Decklin Foster

%
[Om åtgärder för att förhindra fusk i skalvet]Jag menar, så länge jag kan göra mina raketgevär ser ut som en stor Twinkie,Jag skulle bli glad ;)
		-- Qeyser <keyser@jhu.edu>

%
<Knghtbrd> r0bert: kort sagt, vi flyttar flera saker klienten           för närvarande är ansvarig för att berätta servern i saker som           serverkontroller för sig själv<Knghtbrd> Om Neo säger "Det finns ingen sked", The Matrix kommer att säga "Oh ja           Det finns --- inget fusk! "<Hollis> Men han vet kung fu ...<Knghtbrd> Visst han gör, men jag har ett raketgevär.
		-- Qeyser <keyser@jhu.edu>

%
* Kvicksilver lugnt bort XT-Ream arm ..* Kvicksilver fortsätter sedan att slå XT-Ream med XT-Ream arm.<Knghtbrd> wow, är allt detta skalvet hacking gör Mercury våldsam här* Mao är glad skalvet smedjan projektet är i goda händer
		-- Qeyser <keyser@jhu.edu>

%
<Knghtbrd> CVS / Inlägg hade linjen jag behövde "ändra"<Mercury> Knghtbrd: Var på väg att nämna ett sådant .. <G><Mercury> Knghtbrd: Nu redo att begå?<Knghtbrd> önska mig lycka<Knghtbrd> Mercury: det begås<Knghtbrd> Mercury: och efter allt detta, jag skulle vara alltför.
		-- Qeyser <keyser@jhu.edu>

%
* Knghtbrd korsar tårna<Knghtbrd> (om jag korsade mina fingrar skulle det vara svårt att skriva)
		-- Qeyser <keyser@jhu.edu>

%
<Doogie> finns det en dålig sak om att ha en mobiltelefon.<Doogie> Jag kan nås när som helst. : |<Wmono> det är därför jag lämnar min bort hela tiden. ;>
		-- Qeyser <keyser@jhu.edu>

%
<Palisade> hur ska vi uttala '00 eller '01 eller '02 och så vidare?<Deek> Säg adjö till nittiotalet, säga hej till naughties. :)
		-- Qeyser <keyser@jhu.edu>

%
<Deek> Om användaren pekar pistolen mot hans fot och drar avtryckaren, det       är vår uppgift att se till att kulan får där det är tänkt att.
		-- Qeyser <keyser@jhu.edu>

%
<Mercury> Varnas, jag har ett tangentbord jag kan använda för att slå loser huvuden          i, och sedan fortsätta att använda ... (=:]<Deek> Mercury: Åh, en IBM. :)
		-- Qeyser <keyser@jhu.edu>

%
<Palisade> knght, sheesh, du klistrar mina ord ur sitt sammanhang i           #debian eller något?<Palisaden>;)<Knghtbrd> Nej, men jag skulle nog vara;><Palisade> d'oh!
		-- Qeyser <keyser@jhu.edu>

%
<Cas> Mercury: gpm är inte en mycket bra webbläsare. fixa det.
		-- Qeyser <keyser@jhu.edu>

%
<Cas> väl det ya gå. säga något dumt i irc och ha det      förevigade för alltid i någons .sig fil
		-- Qeyser <keyser@jhu.edu>

%
Microsoft är en korsning mellan Borg och Ferengi. Tyvärr,de använder Borg att göra sin marknadsföring och Ferengi att göra sittprogrammering.
		-- Simon Slavin

%
Jag skulle hellre tillbringar 10 timmar att läsa någon annans källkod än 10minuter lyssnar på musak väntar för teknisk support som inte är det.
		-- Dr. Greg Wettstein, Roger Maris Cancer Center

%
Var tror du att du kommer idag?
		-- Dr. Greg Wettstein, Roger Maris Cancer Center

%
Jag hade hört alla typer av dysterhet och doom prognoser för Y2K, så jag trodde jag skulle lyssna några av de råd som experterna har gett: Fyll upp bilens bensintank, fylla på konserver, fylla badkaret med vatten, och så vidare.Jag antar att jag inte var helt vaken när jag avslutat mina förberedelser i slutet av förranatt. I morse hittade jag kökshyllorna indränkt i bensin, vatteni bilens bensintank, och min badkar fyllt med vita bönor.
		-- Dan Pearl in a message to rec.humor.funny

%
<Tarzan> Hej har du faller av din pirch eller något?<Knghtbrd> mig? heh.
		-- Dan Pearl in a message to rec.humor.funny

%
<Espy> du bakat<Knghtbrd> Espy: endast hälften så
		-- Dan Pearl in a message to rec.humor.funny

%
<Darkangel> jag i allmänhet inte använda något som har "experimentell" och            "Varning" klistras över det<Darkangel> nej, jag är inte så dum ... hehe<Knghtbrd> ...* Darkangel anser att hämta den senaste instabil kärna
		-- Dan Pearl in a message to rec.humor.funny

%
<Wichert> solaris är BSD, så det borde fungera* Espy tar Wicherts crack pipe bort
		-- Dan Pearl in a message to rec.humor.funny

%
<Knghtbrd> Det är synd mest gamla Unix visade sig Y2K kompatibel<Knghtbrd> eftersom det innebär att människor kommer fortfarande att köra dem i 30 år           = p<Knghtbrd> det skulle ha varit så mycket trevligare om y2k effektivt dödade av           HPUX, aix, SunOS, etc;><Espy> Knghtbrd: Sedan när är PH-UX, värk och solartus "gamla"?
		-- Dan Pearl in a message to rec.humor.funny

%
* Gxam undrar om alla dessa globals verkligen är nödvändiga<Knghtbrd> flesta av dem just nu ja<Knghtbrd> vi verkligen behöver för att rensa upp dem vid något tillfälle<Knghtbrd> gxam: de globals kommer att behöva gå bort som vi vandrar mot           modularitet och galenskap (dvs libtool)
		-- Dan Pearl in a message to rec.humor.funny

%
<Raptor> Adamel, jag tror koden du fast av mina fungerade inte<Raptor> Jag får inte ha begått arbetskoden<Knghtbrd> raptor: som det är första gången som någonsin har hänt = p
		-- Dan Pearl in a message to rec.humor.funny

%
<Mercury> Knghtbrd: Använda -3dfx eller -svga?<Knghtbrd> Kvicksilver kommer att göra något förnuftigt med det<Knghtbrd> Mercury: båda --- SVGA sig11 s, -3dfx sig4 s<Knghtbrd> Mercury: det är inte bra rätt? ;>
		-- Dan Pearl in a message to rec.humor.funny

%
<Knghtbrd> Lita på oss, vi vet vad vi gör ... Vi kanske inte har någon aning om hur           vi gör det, men vi vet vad vi gör.
		-- Dan Pearl in a message to rec.humor.funny

%
<Mercury> <CJ | Bizkit-0-> jag kan ladda upp till Linux-server tho<Mercury> <CJ | Bizkit-0-> jag fick ett skal konto på en<Mercury> <Mercury> Vad det igång?<Mercury> <CJ | Bizkit-0-> umm<Mercury> <CJ | Bizkit-0-> apache jag tror<Mercury> Hjälp, snälla hjälp ..* Omni skrattar
		-- Dan Pearl in a message to rec.humor.funny

%
<Jt> bör ett fel markeras kritisk om det bara påverkar en båge?<James-workaway> jt: rc för den båge kanske, men dessa slags båge                 specifika buggar är sällsynta ...<Jt> inte när det är på grund av ett fel i gcc<Doogie> JT: få GCC bort från den båge. :)
		-- Dan Pearl in a message to rec.humor.funny

%
<Edlin> LWE?<Edlin> Linux W ?? E ??<Ser> kommer eatyou<JHM> World Expo?<Edlin> jag ser
		-- Dan Pearl in a message to rec.humor.funny

%
"Nominell avgift". Vad en ful mening. Det är en av de saker sominnebär att om du måste fråga, kan du inte råd med det.
		-- Linus Torvalds

%
<Deek> du GPL dina läxor? :)<Knghtbrd> yah = D<Knghtbrd> Alla har rätt att använda eller ändra min läxa, men om de           distribuera förändringar de måste inkludera hela maskinläsbar           källkod;>
		-- Linus Torvalds

%
* Knghtbrd är varje dag mer övertygad om att de flesta C ++ kodare vet inte vad           fan de gör, vilket är anledningen till C ++ har en så dålig rap<CULus> kb: Mest C kodare vet inte vad de gör, bara det gör det        lättare att dölja: P<CULus> se till exempel, proftpd: P
		-- Linus Torvalds

%
<CULus> Och inte få mig började perl!<CULus>:><Shaleh> perl är bortom ont<Jim> du inte vet perl ännu?<Netgod> gotta love språk utan definierbara syntax
		-- Linus Torvalds

%
<Doogie> cat / dev / random | perl?<Shaleh> doogie: det är också ett giltigt sendmail.cf<Doogie> :)* Knghtbrd händer Doogie en meningslös användning-av-katt award* Shaleh vill prova men är rädd
		-- Linus Torvalds

%
<Dhd> perl </ dev / bdsm<Knghtbrd> du har en / dev / bdsm?<Dhd> säker, det är en pseudosadomasochistic slumptalsgenerator
		-- Linus Torvalds

%
<Kysh_> Joey: Jag är på det just nu .. 3 1.3GB skivor, 128M RAM, dubbla 50 Mhz        (Upp till quad 250MHz)<Kysh_> Fångsten är att det drar 110v på cirka 12A 8><CULus> 12A!<CULus> Okej, är min spis 3000W, är denna sol 1320W<CULus> Ser du en PROBLEM HÄR<Calc> en 1320W sol, är det som en hårtork :)
		-- Linus Torvalds

%
* Joeyh_ kör ps och ser 10 rader awk kod* Joeyh_ ryggar i skräck
		-- Linus Torvalds

%
<Knghtbrd> joeyh: Jag var nere sedan förmiddagen igår och PacBell sade           i morse att AT & T var att skylla och nästan alla av staten           var ned<Rcw> vet inte varför folk insisterar på internet kan överleva en kärnvapenkatastrof      när den inte kan överleva en traktorgrävare
		-- Linus Torvalds

%
Detta meddelande skrevs med VI! (Inte att någon i världen bryr sig)
		-- seen on an old message from an anon.penet.fi address

%
återställning anslutning av någon idiot med en traktorgrävare
		-- seen on an old message from an anon.penet.fi address

%
5 februari 13:27:01 treenighet lp0 i brand        - Linux-kärnan, varna mig att det fanns någon okänd           problem med min skrivare (dvs var det slut på bläck)
		-- seen on an old message from an anon.penet.fi address

%
Ju mindre du vet om datorer ju mer du vill Microsoft!        - Microsoft annonskampanj, circa 1996(Bevis att Microsofts reklam _isn't_ oärlig!)
		-- seen on an old message from an anon.penet.fi address

%
Göra ett lysande beslut och en hel massa mediokra sådana är inte såbra som att göra en hel del i allmänhet smarta beslut helahela processen.
		-- John Carmack

%
Det är vanligtvis inte kostnadseffektivt tid klokt att gå göra det. Men om något ärverkligen pissing dig, du bara gå hitta koden och fixa det och det ärväldigt coolt.
		-- John Carmack, on the advantages of open source

%
<Calc> ja det låter bra för RE'ing USB<Calc> Jag har en värdelös 3com USB-kamera här :(<Knghtbrd> calc: 3Com kan få dig arresterad för brott mot lagar som           inte existerar "till oktober;><Beräknat> knghtbrd: Jag kommer att dölja :)<Knghtbrd> ... motstånd gripandet också va?<Beräknat> knghtbrd: nej jag kommer att dölja innan jag få tjänstgjorde
		-- John Carmack, on the advantages of open source

%
<Mercury> Vid den tidpunkten kommer det att sammanställa, men segfault, som det ska ..
		-- John Carmack, on the advantages of open source

%
* Knghtbrd är alltför frestad att .sig hela denna diskussion ...
		-- John Carmack, on the advantages of open source

%
Den Unixverse slutar tis, 19 Jan 2038 03:14:07 0000
		-- John Carmack, on the advantages of open source

%
<Taniwha> Knghtbrd: vi bör göra ett skalv episod: knä djupt i koden ":          du springa runt skjuta på fel :)<Knghtbrd> Taniwha: Jag ska förmedla idén till OpenQuartz;>
		-- John Carmack, on the advantages of open source

%
<Taniwha> jag skulle lösa en Windows-tangenten problem med fdisk :)
		-- John Carmack, on the advantages of open source

%
<Endy> knghtbrd: QW s netcode gör konstiga saker till mig. : P<Knghtbrd> Detta är ovanligt? ;><Endy> Inte riktigt. : P
		-- John Carmack, on the advantages of open source

%
<Knghtbrd> rcw: Åh yay --- Jag har inte varit inblandad i en bra gräl in på           minst ... 5 minuter!
		-- John Carmack, on the advantages of open source

%
<Manoj> shaleh: Jag är inte, trots din förstått Gud
		-- John Carmack, on the advantages of open source

%
<SlayR> Jag har precis köpt MS Office 2000 för endast $ 20 !!!<Knghtbrd> du fick rippat;><SlayR> jag vet;)
		-- John Carmack, on the advantages of open source

%
<Knghtbrd> det är 06:00. Jag har varit upp 24 timmar<Knghtbrd> Vakna mig upp och risken liv och lem.* Knghtbrd &; sova<Tv> Okej alla, vi vänta 10 minuter och sedan börja översvämningar Knghtbrd     med ^ G. Någon hacka rot och katt / dev / urandom> / dev / dsp.
		-- John Carmack, on the advantages of open source

%
*** Knghtbrd är nu känd som SirKewLDooD*** Kvicksilver sparkas SirKewlDooD från #quakeforge (* FÖRSÖK *)
		-- John Carmack, on the advantages of open source

%
<Mercury> Knghtbrd: Jag skulle gärna vilja se stöd för XOR hårkors ..<Knghtbrd> Mercury: du är på kvacksalvare.<Mercury> Knghtbrd: Du är återförsäljaren ... <G>*** Knghtbrd är nu känd som QuackDealer
		-- John Carmack, on the advantages of open source

%
* Torris kan inte koda sin väg ut ur en papperspåse<Coderjoe> torris: int main () {ExitPaperBag (); tillbaka 0; }<Knghtbrd> Är det hur det är gjort då? * Tar anteckningar *
		-- John Carmack, on the advantages of open source

%
<Knghtbrd> eek, inte en annan ...<Knghtbrd> Verkar någonsin utvecklare och deras mor har nu en slumpmässig           signatur använder irc citat ...<Knghtbrd> vad har jag började här ??
		-- John Carmack, on the advantages of open source

%
* Ser använder knghtbrd kommentarer som hans signatur<Knghtbrd> ser: så fort jag skrivit dem insåg jag att jag skulle bättre klippa dem           själv innan någon annan gjorde;>
		-- John Carmack, on the advantages of open source

%
* Omnic tittar på sin 33,6 länk och sedan tittar på Joy* Kvicksilver kelar hans kabelmodem .. (=:]
		-- John Carmack, on the advantages of open source

%
Visst, Win95 utseende var inte allt det nya antingen - Apple försökte att stämmaMicrosoft för att kopiera Macintosh UI / papperskorgen, tills Microsoftpåpekade att Apple fick många av sina Mac idéer (inklusive papperskorgenikon) från Xerox ParcPlace. Xerox förmodligen fortfarande undrar varföralla är intresserade av sina soptunnor.
		-- Danny Thorpe, Borland Delphi R&R

%
<Knghtbrd> är det ett tecken på psykisk sjukdom att vandra planlöst genom           börja karta, samla in din Thunderbolt, hoppa i poolen, och GIB           dig med det bara för att se huvudet buouce när det fallergenom botten av poolen? =><Knghtbrd> "Du vet att du är en Quake missbrukare när ..."
		-- Danny Thorpe, Borland Delphi R&R

%
<Zoid> Jag tror fortfarande att ni är nötter sammanslagning Q och QW. : P<Knghtbrd> Naturligtvis är vi nötter. Även John sa det. =><Taniwha> Zoid: vi är nötter, men vi är produktiva nötter :)
		-- Danny Thorpe, Borland Delphi R&R

%
<Taniwha> Zoid: vi är nötter, men vi är produktiva nötter :)* Taniwha undrar vad produktiva nötter smakar
		-- Danny Thorpe, Borland Delphi R&R

%
<Endy> Taniwha: Citat material :)<Taniwha> Endy: :)<Knghtbrd> Endy: Jag har redan klippt det
		-- Danny Thorpe, Borland Delphi R&R

%
<Endy> Faktiskt, jag tror att jag ska vänta på potatis att slutföras före       installera debian.<Endy> Det borde vara snart, jag hoppas. :)<Knghtbrd> Endy: Du vet uppenbarligen mycket lite om Debian.
		-- Danny Thorpe, Borland Delphi R&R

%
Ingenting är ett problem när du felsöka koden.
		-- John Carmack

%
<Overfiend> Unix sätt - allt är en fil<Overfiend> Linux vägen - allt är ett filsystem :)
		-- John Carmack

%
<Devkev> Ja jag såg blixten pistol och där ni skulle, tänkande         du skulle sparka några ass :)<Devkev> insåg att det skulle vara din egen :)
		-- John Carmack

%
"Annars, tala med en läkare om att ta bort huvudet frånröv, tror jag att det skulle vara till fördel för alla inblandade. "
		-- Zephaniah E. Hull, flaming someone on a mailing list

%
Tagline, är det!
		-- Zephaniah E. Hull, flaming someone on a mailing list

%
Jag tränar en fin punkt etik. Det är acceptabelt att skjuta tillbaka.Det är inte acceptabelt att skjuta först.
		-- Zed Pobre

%
<Coderjoe> gib, perl?<Gib> methinks perl är programmerarens schweiziska armé Chainsaw
		-- Zed Pobre

%
<Endy> Taniwha: Har du testat den här en? :)<Taniwha> Endy: naturligtvis inte
		-- Zed Pobre

%
Det är det roligaste jag någonsin har hört och jag kommer _inte_ tolerera det.
		-- DyerMaker, 17 March 2000 MegaPhone radio show

%
Det är inte? Menar du att du bör tillåta människor (andra än WilliamWallace) att skjuta blixtar från sin åsna?
		-- Seth Galbraith

%
<Mercury> Du behöver inte vara galen för att vara en medlem av projektet, men          du kommer att bli .. <=:]
		-- Seth Galbraith

%
* Endy måste rådgöra kaffe: P<Endy> kaffe bot personen, inte kaffe drycken :)<Knghtbrd> samråd drycken kan hjälpa också =>
		-- Seth Galbraith

%
<Mongoose> knghtbrd: och de ödmjuka skall ärva K-Mart
		-- Seth Galbraith

%
<Knghtbrd> "Java för COBOL programmerare"<Knghtbrd> som skriver dessa saker?<raptor> folk på crack<raptor> och COBOL programmerare<Raptor> :)<Knghtbrd> som är överflödig.
		-- Seth Galbraith

%
<Evilkalla> heh, jag tog aldrig en kodnings klass<Evilkalla> eller en grafisk klass<Evilkalla> eller en mjukvarudesign klass<Vegan> och det visar: P
		-- Seth Galbraith

%
* The_Answer_MD kastar spaghetti på alla* Taniwha äter spaghetti* Coderjoe kastar runt några köttbullar* Knghtbrd får osten* Taniwha griper en röd
		-- Seth Galbraith

%
<Theoddone33> Vad är detta meddelande på skärmen,<Theoddone33> så blå, så blå, vad kan det betyda?<Theoddone33> Kan ni, skulle du trycker på Radera<Theoddone33> Ctrl och Alt och sedan upprepa.
		-- Seth Galbraith

%
<Gorgo> vad du får när någon sprickor din debian maskin?<Gorgo> potatismos ...
		-- Seth Galbraith

%
<Aj> komma på<Aj> det är en pico-klon<Aj> det * betydde * att vara irriterande
		-- Seth Galbraith

%
<Espy> Jag åberopar Espy lag, som säger att ni suger: P
		-- Seth Galbraith

%
<Overfiend> cULus: vill avbryta mig för det? :)<CULus> Overfiend: Gå skadligt knäcka några klipper och vi pratar<Overfiend> cULus: Fan, måste det vara skadlig?<CULus> Overfiend: Tyvärr ja
		-- Seth Galbraith

%
<Knghtbrd> 2fort5 suger nog att ha sin egen gravitation ...
		-- Seth Galbraith

%
* Kosmiska partiklar önskar att han hade några strippor här ....<Kosmiska partiklar> fela, Avisoleringstänger
		-- Seth Galbraith

%
<Wildthing> ok killar .. så whens nästa begå: PP<Taniwha> när de kommer att få mig
		-- Seth Galbraith

%
<Mdorman> Jag är en gnuer personen själv. Det är en redaktör! Det är en floorwax!          Det är en dessert toppning!
		-- Seth Galbraith

%
<Tausq> F. Vad är skillnaden mellan Batman och Bill Gates?<Tausq> A. När Batman kämpade Penguin, han vann.
		-- Seth Galbraith

%
Vid något tillfälle, bitar måste gå in paket och routrar måste görabeslut om dem. Förändringar på den nivån är vad jag vill höra om, intestrategiska företag relationer.
		-- John Carmack

%
Vi avvisar: kungar, presidenter, och rösta.Vi tror på: grov konsensus och arbetskoden.
		-- Dave Clark

%
<Knghtbrd> QF kommer att få zipfile stöd idag<Coderjoe> heh ... InfoZip?<Knghtbrd> Har jag tur ja<Deek> knghtbrd: Du skojar, va? ;)* Deek tar bort Knghtbrd s crack pipe. ;)
		-- Dave Clark

%
<Deek> ändra alla cvar-> värde = X att använda Cvar_Set ()<Theoddone33> som inte skedde i oldtree<Deek> Egentligen gjorde det.<Knghtbrd> ja - två veckor senare.
		-- Dave Clark

%
=== Detta brev är Honor System Virus ====Om du kör en Macintosh, OS / 2, Unix, ellerLinux-dator, vänligen slumpmässigt ta bortflera filer från hårddisken ochvidarebefordra detta meddelande till alla du känner.==============================================
		-- Dave Clark

%
* Genväg vill få i en av knghtbrd s sigs en av dessa dagar.
		-- Dave Clark

%
<Dr ^ Nick> SGI_Multitexture är dålig voodoo nu<Dr ^ Nick> ARB är bra voodoo<Witten> nej, voodoo rusa dålig voodoo :)
		-- Dave Clark

%
99 små buggar i koden, 99 buggar i koden,        fixa en bugg, kompilera det igen ...        101 små buggar i koden ....
		-- Dave Clark

%
Hmm ... Vilket skulle göra ett bättre jobb på att köra fysiker galen? Resasnabbare än ljuset, eller en flyttals booleskt värde?
		-- Michael Mol

%
<Beräknat> knghtbrd: gnome 2.0 kommer vara ute i ett par månader, inte säker på hur det       kommer att jämföra med kde 2,0 men<Knghtbrd> calc: Lika uppsvälld, precis som buggig, och varje Gnome 2 app       kommer att bero på 30 bibliotek.<Slimer> knghtbrd: så vilka förändringar från 1,0?
		-- Michael Mol

%
<Ze0> så, hur är allt i världen av Quack?<LordHavoc> Precis Ducky<Ze0> utmärkt, stekt anka är mighty fine välsmakande.
		-- Michael Mol

%
<FrikaC> Jag borde starta ...<FrikaC> OK brb<FrikaC> Så, vad isär formen undvika virii, minnesläckor och frodas         krascha gör Linux reallhy erbjuda :)<LordHavoc> tillförlitlig multitasking?
		-- Michael Mol

%
<Tausq> if (cb) ((CB> obj) -> * (CB> ui_func)) ();<Knghtbrd> tausq: Vem fan skrev det?<Tausq> mig :)* Knghtbrd flogs tausq
		-- Michael Mol

%
<Knghtbrd> glDisable (GL_BUGS);<Endy> heh<Endy> Är det i 1.2? :)
		-- Michael Mol

%
<Mercury> knghtbrd: Eww, hitta ett bättre namn, suger filmen .. <G><Knghtbrd> Mercury: Motorn är bättre än filmen
		-- Michael Mol

%
<LackOfKan> Vad är "bots"?< `` Erik> RSG är en bot, inte en människa, inte en mänsklig användbar klient, bara en bot.< `` Erik> ungefär samma som ett skalv bot, utom irc bots är (oftast)         byggd för att hjälpa, inte skjuta din röv full av hål
		-- Michael Mol

%
if (mig = dig!) // FIXME: förmodligen alltid sant, ta bort?    för (n = 0; n <who_knows_what; n ++) {        answer = doSomething (withthis [n]);        if (svar == foobar) {            GetLost (n);            ha sönder;        }    }
		-- Michael Mol

%
<Knghtbrd> Yorick: inga problem med indexerade färgpaletter för bilder, som           länge du kan plocka paletten<Yorick> Uppenbarligen människor skapar skalvet var färgblind, men det         betyder inte att du måste vara
		-- Michael Mol

%
<cesarb> Fan, varje gång jag leka, QF-client-x11 lås hårt<Zoid> inte dö?<Knghtbrd> bra incitament.
		-- Michael Mol

%
Varför är det att alla de instrument som söker intelligent liv iuniversum är pekade bort från jorden?
		-- Michael Mol

%
<Rebelpacket> Hej, snabb fråga, finns det något sätt att påskynda              prestanda uquake-x11?<Deek> rebelpacket: Om du vill påskynda den, kasta det svårare.
		-- Michael Mol

%
<Netgod> du vet<Netgod> dess verkligen sorgligt när InterNIC själv inte kan konfigurera DNS         servrar rät<Netgod> det bara blir inte mer patetiskt än
		-- Michael Mol

%
<Knghtbrd> Även med overbrights är Quake färgpalett full av tråkig,           platta färger<LordHavoc> knghtbrd: skalvet palett är mycket levande om du inte använder gamma            korrektion<LordHavoc> väl egentligen håller jag, det är långt ifrån lika levande som Unreal<Deek> Q3 å andra sidan ... NEON.<LordHavoc> Q3 är bara löjligt<Deek> Q3 tar medeltida kyrkfängelsehåla och lägger det i Vegas.
		-- Michael Mol

%
"Jag har ett ben att plocka, och några att bryta."
		-- Anonymous

%
Z.O.I.D .: Zombie Optimerad för Infiltration och Destruction
		-- Anonymous

%
<Deek> Ja, är Amerika ett land beroende på hur förbannad-off en grupp beskattas       människor kan få.<Deek> Vi finns som ett land eftersom vi är billig.
		-- Anonymous

%
<Oskuro> Overfiend: många fläckar på toppen av 4.0.1 redan?<Overfiend> Oskuro: ett fåtal<Overfiend> endast 152 meg
		-- Anonymous

%
<Joeyh> oh my, är det en UPP P III.<Doogie> dos den.* Joeyh löper dselect<Overfiend> som borde vara tillräckligt :)
		-- Anonymous

%
<Barneyfu> knghtbrd: skit, gör SDL säker DGA en jävla massa lättare för           inte det? :)<Knghtbrd> barneyfu: vad DGA?<Barneyfu> mus DGA<Knghtbrd> barneyfu: (inte att svara på din fråga?)<Barneyfu> hahahahaha YEAH! :)
		-- Anonymous

%
<Deek> "En bra programmerare kan skriva FORTRAN på alla språk."<Deek> knghtbrd har visat att du kan skriva C ++ på något språk också.       <Grin><Mercury> Vi håller considdering om vi skulle ge honom eller pris, eller          döda honom..<Mercury> (Naturligtvis, med alla rättigheter, innebär det att vi skulle ge honom          pris, och sedan döda honom .. <G>)
		-- Anonymous

%
En omstörtande är någon som kan ut-argumentera för sin regering.
		-- Anonymous

%
Vi måste veta, vi kommer att veta.
		-- David Hilbert

%
<Knghtbrd> Internet censur. Eftersom dina barn måste vara           skyddad från nakna kvinnor, medicinska procedurer, diversekulturer och våldsamma videospel.<Knghtbrd> (men information om att bygga bomber, stjäla kabel, och           tillverka läkemedel är okej ...)
		-- David Hilbert

%
En vän till mig har en streckkod på armen.Han ringer upp som en $ 0,35 pack JuicyFruit.
		-- Seen on Slashdot

%
<NullC> Jag gillar fröet kod för att beräkna maskeringskurvor.<NullC> Jag har aldrig sett kod som gjorde att vill dricka innan ...
		-- Seen on Slashdot

%
$ Du = ny DIG;tuta () om $ dig-> love (perl)
		-- Seen on Slashdot

%
<Cj> nej! problem i M $ programvara?<Cj> "Grundligt bugtested"* Dabb flinar.<LordHavoc> skriva om det såsom "Grundligt buginfested '
		-- Seen on Slashdot

%
<Doogie> dpkg har buggar? aldrig!
		-- Seen on Slashdot

%
"Debian: inga hattar eller reptiler harmed i danandet av denna fördelning =. "
		-- Paul Slootman

%
* Athener kallar Amnesty International House of Pancakes
		-- Paul Slootman

%
<Elmo> oren fela, admin laget kontrollerar inte arkivet, det är       ftp cabal<Elmo> få dina cabals rätt, fan det :-P
		-- Paul Slootman

%
<Benc> kosmiska partiklar: du fylla mig<Benc> err ...<Kosmiska partiklar> heh* Benc går tillbaka till kodning* Elmo tittar på Benc<Elmo> något som vi bör veta om dig och kosmiska partiklar, Ben? :)
		-- Paul Slootman

%
Ändra det sociala kontraktet? BWAHAHAHAHAHAHAHAHAHAHAHA.
		-- Branden Robinson

%
<Knghtbrd> Program mottagna signalen SIGSEGV, Segmente fel.<Knghtbrd> 0x40095fb0 i memchr () från /lib/libc.so.6<Knghtbrd> (GDB) bt<Knghtbrd> # 0 0x40095fb0 i memchr () från /lib/libc.so.6<Knghtbrd> # 1 0x0 i ?? ()<Knghtbrd> Jo det är verkligen till hjälp* Knghtbrd handlar gdb för en trevlig ouija ombord - det hjälper mer
		-- Branden Robinson

%
Alla goda idéer ser ut som dåliga idéer till dem som är förlorare.
		-- Dilbert

%
RFC 882 sätter pricken i .com, inte Sun Microsystems
		-- Seen on Slashdot

%
* Joeyh_ undrar om Linux är tänkt att låsa upp när du frågar 100  processer för katt hela cd-enheten
		-- Seen on Slashdot

%
<Pretzelgod> knghtbrd: Quake bör stödja xray vision, dammit<Knghtbrd> pretzelgod: ftp://ftp.cdrom.com/pub/quake/partial_conversions/           xrated / i_am_old_enough_to_look_at_this<Knghtbrd> ... du frågade ...<Kosmiska partiklar> haha, är att en riktig katalog
		-- Seen on Slashdot

%
<Knghtbrd> I smyga Bun<Knghtbrd> hjälpa mig för ATT kvacksalvare<Venom> kb: vad fan pratar du om?<Knghtbrd> bwahahaha .. Det är en lång historia.
		-- Seen on Slashdot

%
<WildCode> Kvicksilver, inte felsökning X lite som att hitta perfekt           Bugffri koden i fönster ??<Mercury> WildCode: Debugging X är som att försöka köra en rak linje          genom en labyrint.<Mercury> Du behöver bara böja rumtiden så att hörnen flytta runt          dig och du kommer inte ha några problem. (=:]
		-- Seen on Slashdot

%
<Miguel> 'Du har varit prenumerationen på hög energi personlig         skyddsanordningar e-postlista "<Miguel> Jag minns att komma in sändlistan inte
		-- Seen on Slashdot

%
<Myt> Jag får en förbindelse vägrade när du ansluter till port 25, någon       vet var fan stocken är?<Aj> Myt: /var/log/damn.log?* Aj undrar vad som skulle se ut<Aj> 18 december 05:32:30 Blåe smtpd [123]: Fan allt TO HELL !!
		-- Seen on Slashdot

%
* Vessla undrar hur dum man måste vara att spam alt.anonymous.messages<Knghtbrd> vessla: ungefär hälften så dum som man måste vara för att skörda den.
		-- Seen on Slashdot

%
* Wolfie funderar hur många Debian det tar att skruva i en glödlampa<Viiru> wolfie: Någonstans runt 600? En skruv är glödlampan, och resten        flamma honom för att göra fel.<Del> wolfie: är lampan fri programvara?<Tv> Kan vi rösta om att skruva eller inte?
		-- Seen on Slashdot

%
<Culus_> Vi hoppas också att släppa en version av Linux där skalet är         ersättas av perl i hög grad. Lägga till att det finns en         Några av oss som vill se en ren perl plattform .. Perlos :)* Culus_ ser på i skräck<Mstone> Culus_: på sidan upp du kan skriva fan nära någonting på         kommandotolken :)
		-- Seen on Slashdot

%
<Mercury> LordHavoc: Anledningen till GL har övertrassera beror på att det är endast          användning av halva det system som de utformats för vis.<Mercury> LordHavoc: Skytte själv i foten.* Dabb tittar på alla dessa kulhål i skorna - jävla, massor :)
		-- Seen on Slashdot

%
<Dabb> hehe, jag hatar verkligen felrapporter som är som ringer brand       avdelning och säger: "Det är eld hit, kom" :)<Dabb> (och hänga upp)* Dabb dödar dussin felrapporter.
		-- Seen on Slashdot

%
<Xtifr> wow, jag tror att jag bara använde libtool för att lösa ett problem - någon        hjälp mig! :><Luca> xtifr, steg bort från tangentbordet
		-- Seen on Slashdot

%
<Mao> varför de insisterar på ading -Werror ...<Misty-chan> Mesa inte skulle kompilera ur lådan om det gjordes av dig             guys;)<Knghtbrd> Uh, Mesa INTE sammanställa ur lådan för det mesta.
		-- Seen on Slashdot

%
<Deek> nopcode: Nej, det är inte. Win32 saknar motsvarande fork ().<Knghtbrd> Deek: windoze är inte avsedd för personer som ska ha tillgång till           vassa föremål, varför ingen gaffel ()<Knghtbrd> istället, måste du lita på sked ()
		-- Seen on Slashdot

%
<Knghtbrd> Detta typsnitt börjar komma ut mycket snyggt<Stu> Knghtbrd: Åh kära, du hacka upp en annan skalvet teckensnitt i VI? :)
		-- Seen on Slashdot

%
<Pv2b> oh, förutom, vad det bästa tillvägagångssättet om jag vill göra en Quake       nivå som utformats från en befintlig byggnad?<Knghtbrd> Få en planlösning av Brian kontor? =)<Pv2b> Knghtbrd: im med tanke på min skola.<Knghtbrd> Oh great<Knghtbrd> Det är allt vi behöver
		-- Seen on Slashdot

%
<Knghtbrd> Windoze Cement: Nu med CrackGuard (TM)! Aldrig oroa           fula sprickor i Windoze cement igen! CrackGuard (TM) ärså kraftfull att det hela kommer att falla sönder innan den kommerspricka. Beställ din $ 200 uppgradering idag!
		-- Seen on Slashdot

%
<Doogie> cULus: min bugg med OpenSSH verkar vara fast i 2.5.2, men         befälhavaren körs 2.3.0<CULus> Inte ens starta<Doogie> Jag gjorde bara.<CULus> Ni kommer att köra mig att bygga en stor gigantisk robot och        förstöra alla Texas, är inte du?
		-- Seen on Slashdot

%
<Shader> vad fel med rjing?<Rhamphoryncus> det är lame: P<Rhamphoryncus> Det bör inte vara möjligt<Rhamphoryncus> prejar en granat upp din röv och använder den som raket                drivmedel bör inte vara en livskraftig teknik: P
		-- Seen on Slashdot

%
 * Motsvarande kod är tillgänglig från RSA Data Security, Inc. * Denna kod har testats mot det, och motsvarar, * Förutom att du inte behöver omfatta två sidor av legalese * Med varje kopia.
		-- public domain MD5 source

%
* Knghtbrd är borta - zzz - meddelanden kommer att snappas som våta handdukar på alla  av de människor som har stulit varumärket knghtbrd frånvaromeddelande<Coderjoe> ack* Coderjoe förbereder sig för att försvara sig från våta meddelanden
		-- public domain MD5 source

%
Underskatta aldrig kraften av någon med källkod, en textredigerare,och viljan att helt slang deras system.
		-- Rob Landley <telomerase@yahoo.com>

%
"Så kommer Andover partiet har en kontant bar?""Nej, det är gratis öl.""Uh-oh, Stallman kommer att bli förbannad ..."
		-- overheard at the Bazaar, 1999

%
<Addi> Alter.net verkar ha ersatt en av dess router med zucchini.
		-- overheard at the Bazaar, 1999

%
<Mercury> Någon fixa det.<Förtvivlan> begåtts<Knghtbrd> förtvivlan: Mercury?<Förtvivlan> Knghtbrd: han är trött, gjorde ett misstag, ville att någon skulle ångra det.<Knghtbrd> förtvivlan: så att du hade honom begått?<Förtvivlan> Knghtbrd: ja, tillägnad ändå.
		-- overheard at the Bazaar, 1999

%
<Taniwha> Knghtbrd: det är inte svälla om det används<Knghtbrd> Taniwha: Hur förklarar ni windoze då?<Taniwha> Knghtbrd: det mesta används endast som ballast för att se till att din          hårddisk är full<Knghtbrd> Taniwha: ballast ... Är inte det vad som gör subs sjunka till           botten av havet?<Knghtbrd> Taniwha: som skulle förklara varför winboxes alltid kommer ner.
		-- overheard at the Bazaar, 1999

%
förnya / IN ingen vait / vb .: 1. lämplig tredjepartsteknikgenom köp, imitation eller stöld och integrera den i ende-facto monopol-ställning produkt. 2. För att öka i storlek eller komplexitetmen inte i verktyget; att minska kompatibilitet eller interoperabilitet. 3. Om du villlockout konkurrenter eller att låsa in användarna. 4. För att ta ut mer pengar; tillhöja priserna eller kostnader. 5. För att få vinster från investeringar i andraföretag men inte direkt produkt eller service. 6. För att kväva ellermanipulera en fri marknad; att förlänga monopolrättigheter till nya marknader. 7.Att undgå ansvar för felsteg; att få bort. 8. köplagstiftning, lagstiftare, lagstiftande eller chefer stats. 9.medla alla transaktioner i en global ekonomi; att förskingra; att adjungera makt(statskupp). Jfr förnya, engelsk användning (antonym).
		-- csbruce, in a Slashdot post

%
Det öronbedövande tystnad lärde mig att inte ställa en massa nördar för rådfrån sina flick
		-- csbruce, in a Slashdot post

%
"Vad ska vi göra i kväll, Bill?""Samma sak som vi varje kväll Steve, försök att ta över världen!"
		-- csbruce, in a Slashdot post

%
<Deek> Det påminner mig, vi måste köpa en motorsåg för kontoret. "I       nödfall, krossa glas "
		-- csbruce, in a Slashdot post

%
<Knghtbrd> Han är en ungefär hälften så stor som de andra.<Knghtbrd> Men han har en motorsåg.
		-- csbruce, in a Slashdot post

%
<Deek> "Jag håller mina personliga gpg data i en låst, leder säkert i ett valv       vaktas av arga rednecks och deras dawgs. Inkräktare kommer att vara       kränks, och allt det där ... "
		-- csbruce, in a Slashdot post

%
<Ex Machina> glQuakeIIIRendererMode (GL_TRUE)<Knghtbrd> Ex Machina: är inte den del av förlängningen som ger           glDriverBugs (GL_FALSE); ?<Siigron> Knghtbrd: nej, glDriverBugs () är en del av EXT_help_me.<Siigron> som också innehåller glMakeItWork (GL_PLEASE);
		-- csbruce, in a Slashdot post

%
< `` Erik> 18.446.744.073.709.551.616 är ett stort antal
		-- csbruce, in a Slashdot post

%
<Xavvy> är det verkligen knghtbrd?<Knghtbrd> Nej, jag är en ond SKOJARE!<Knghtbrd> En ond bedragare som gillar HYBRID!<Xavvy> haha<Xavvy> ok, det är honom: P
		-- csbruce, in a Slashdot post

%
<| Regn |> I * love * SWB !!<| Regn |> Eller tryck 5 för att tala med en representitive ..<| Regn |> * 5 *<| Regn |> Du överförs, vänligen håll ...<| Regn |> ...<| Regn |> ...<| Regn |> Tyvärr, detta nummer kan inte slutföras som rings upp.<| Regn |> Kontrollera numret och försök igen.
		-- csbruce, in a Slashdot post

%
<| Regn |> #define struct union / * stort utrymme sparare * /
		-- csbruce, in a Slashdot post

%
<Elric> inga BSD fans?<EvilTypeGuy> Elric: det är svårt att vara en spelare och en BSD fan: p
		-- csbruce, in a Slashdot post

%
<Marticus> Det finns för mycket blod i mitt koffeinsystem.
		-- csbruce, in a Slashdot post

%
<SirDibos> cULus: är du vaken?<CULus> nej
		-- csbruce, in a Slashdot post

%
<WLI> Ja, jag tittade på esd och det såg ut som vilken typ av C-kod som en      ex-JOVIAL / Algol '60 kodare som hade tillbringat de senaste 20 åren studsar      mellan Fortran-IV och Fortran '77 skulle skriva.
		-- csbruce, in a Slashdot post

%
<Olinjära> NET är Microsofts perverterad version av en java nätverks            miljö uglified för Windows-specifik skit
		-- csbruce, in a Slashdot post

%
<Mercury> LordHavoc: Jag är redan galen.<Coderjoe> jävla rakt. eller kurviga, krokiga, eller vad har du
		-- csbruce, in a Slashdot post

%
Unix är mogen OS, Windows är fortfarande i blöjor och de luktar illa.
		-- Rafael Skodlar <raffi@linwin.com>

%
<Midgar> Från alla sterotypes om Aussies, jag räkna ni är         riktigt tuff.<Midgar>; p<Krusto> vi kastar Koalas på dig
		-- Rafael Skodlar <raffi@linwin.com>

%
<| Regn |> * nod * Jag är inte förtjust i att använda smarta värdar, själv<| Regn |> eftersom den bygger på både fjärrvärden och din värd att vara smart<| Regn |> och alltför ofta du missar en av dessa båda mål
		-- Rafael Skodlar <raffi@linwin.com>

%
Sourceforge tillvägagångssätt är att placera alla projekt i några intetsägande"Open source surburbia", där alla husen är likadana, med endastfärger och mindre stilvarianter (vilka byggnadsplan användes somsärskilt hus) tillåts av de restriktiva förbund och lokalazonindelning lagar. Sourceforege är öppen källkod motsvarighet tillindelning i filmen "Edward Scissorhands".
		-- Terry Lambert

%
<Beräknat> Knghtbrd: irc inte kompilera C-kod mycket väl;)
		-- Terry Lambert

%
* | Regn | förbereder sig för polygon soppa<| Regn |> söt barmhärtig skit, fungerar det?* | Regn | svimningar
		-- Terry Lambert

%
"Eftersom det är en självklarhet att Microsoft kommer att vara nedskräpning sin XMLmed pekare till Win32-baserade komponenter, det bästa som kan sägas omdess antagande av XML är att det kommer att göra det lättare för webbläsare ochapplikationer på icke-Windows-plattformar för att förstå vilka delar avdokumentera det måste bortse från. "
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
<Robert> Jag förstår att det finns några rimliga gränser för yttrandefriheten i         Amerika, till exempel jag inte kan skrika Brand i en fullsatt teater.. Men kan jag skrika brand i en teater med bara 5 eller 6 heltidsarbete	 i det ?
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
<AAV> kaffe på fastande mage är ganska nasy<Knghtbrd> AAV: tid att köra till automaten för cheetos<AAV> cheetos? :)
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
<| Regn |> med sane kod, kanske jag kunde räkna ut återgivnings :)<LordHavoc> regn: Jag skulle förmodligen vara en skriva återgivnings<| Regn |> väl, er, eh
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
<| Regn |> Knghtbrd: Låt mig ge dig tillgång till zonfiler<Knghtbrd> oh gudar - du inser jag har aldrig spelat med bind rätt?<| Regn |> uhoh :)
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
<F00Dave> Titta avvisar detta är #OpenGL, inte #GEEKSEX.
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
* TwingyAFK är shopping för 17 "platt* AAV säljer TwingyAFK en bit av plywood
		-- Nicholas Petreley, "Computerworld", 3 September, 2001

%
Är det inte pinsamt när du måste gå till apoteket för vissa"speciella föremål" och när du checkar ut, ser kassören på digsom, "Åh, jag vet vad du gör i kväll ..."Japp, det kassörskan läsa alla tecken ... konserverade kycklingsoppa, Theraflu,Halls, NyQuil de bigass flaskor EGT och grapefruktjuice ... han vissteoch jag visste att jag hade ett datum med teevee och ett duntäcke. awwwja.
		-- Elizabeth Kirkindall

%
Inom vetenskapen det händer ofta att forskare säger, "Du vet att det är en riktigtbra argument; Min ståndpunkt är felaktig, "och sedan de faktiskt ändrasderas sinnen och du hör aldrig den gamla vy från dem igen. de verkligengör det. Det händer inte så ofta som det ska, eftersom forskarna ärmänsklig och förändring är ibland smärtsamt. Men det händer varje dag. Jag kan inteminns förra gången något sådant hände i politik eller religion.
		-- Carl Sagan, 1987 CSICOP keynote address

%
<Knghtbrd> lägga till en GF2 / 3, en betydande hårddisk, och en 15 "platt och           du har en ganska förbannat bärbar maskin.<Coderjoe> en GeForce två tredjedelar?<Knghtbrd> Coderjoe: ja, ett GeForce två tredjedelar, det vill säga något kort från ATI.
		-- Carl Sagan, 1987 CSICOP keynote address

%
<Knghtbrd> Nintendo förklarar GCN populäraste konsolen någonsin<Knghtbrd> Vilka är de skojar?<Mercury> knghtbrd: lager innehavare?
		-- Carl Sagan, 1987 CSICOP keynote address

%
<LordHavoc> majoriteten av windoze konstnärer inte har förmågan att            spara xpm<Mercury> LordHavoc: De har inte anteckningsblock? * G, D & R *
		-- Carl Sagan, 1987 CSICOP keynote address

%
Linux stöder idén om en kommandorad eller ett skal av samma skälatt endast barn läsa böcker med bara bilder i dem. Språk, vare sig detEngelska eller något annat, är det enda verktyg tillräckligt flexibel för att åstadkommaett tillräckligt brett spektrum av uppgifter.
		-- Bill Garrett

%
## Signoff: uppror (razzin "frazzin" motherfu ... dum DirectX ...)
		-- Bill Garrett

%
<Krogoth> Kgnghtbrd: Jag skulle inte kow, jag ser inget behov av en stavningskontroll ännu<Knghtbrd> du sa?
		-- Bill Garrett

%
<Knghtbrd> Jag skulle bättre sätta komprometterande saker i koden: ahfuiovka           ikperoa edfr ade 9 enbuw ejasxleme ka Iena df4mesa<Knghtbrd> Om du kan dekryptera det, du är en bättre cryptographer än jag           am. =)
		-- Bill Garrett

%
<Rcw> liiwi: printk ( "CPU0 eld \ n");
		-- Bill Garrett

%
<Electro> min dator var en gång en av byggstenarna i en stor          pyramid
		-- Bill Garrett

%
OBSERVERA: någon sett röka kommer att antas vara i brand och kommer att vara        summariskt släcka.
		-- Bill Garrett

%
<Markm> c ++: kraften, elegans och enkelhet av en handgranat
		-- Bill Garrett

%
<Knghtbrd> men en sort per flik och ingen per lista är utan tvekan bättre än           O (n + n ** 2) per flik och O (n ** 2) per lista.<Knghtbrd> OMG, någon skjuta mig.<Coderjoe2>?<Knghtbrd> Jag kan inte tro jag bara använt den stora svan ägg för att förklara varför min           sätt är förmodligen bäst i det långa loppet.
		-- Bill Garrett

%
<Hoponpop> mitt program fungerar om jag tar ut buggar.
		-- Bill Garrett

%
<Mercury> Knghtbrd: Hej, har perl effekt grace och elegans av en släde          hammare. (=:]<| Regn |> säkert nåd och elegans, i alla fall
		-- Bill Garrett

%
<DannyS> Hit apan att vinna $ 20 (*)!* Knghtbrd får ut sin klubba.* Knghtbrd växter den ordentligt på DannyS 'huvud.* Knghtbrd tar hans $ 20 nu. = D
		-- Bill Garrett

%
<Gholam> och jag är imponerad<Gholam> win98 lyckats krascha X inifrån VMware.* Gholam applauds.
		-- Bill Garrett

%
"Nvidias drivrutiner för OpenGL är min" gold standard ", och det har varit ganskatag sedan jag har haft att rapportera ett problem för dem, och även deras varumärkenya tillägg fungerar som dokumenterats första gången jag prova dem. När jag harett problem på ett Nvidia, jag antar att det är mitt fel. Med någon annansdrivrutiner, jag antar att det är deras fel. Detta har visat sig korrekt nästanhela tiden."
		-- John Carmack

%
Libtool delade bibliotek portabilitet är endast något mer trovärdigt änevighetsmaskiner. Speciellt på AIX :). "
		-- David Leimbach

%
<Overfiend> detta är den nya Overfiend, predikant kärlek och tolerans
		-- David Leimbach

%
<Hoponpop> skillnaden mellan NetBSD, FreeBSD och OpenBSD, som en           insider är FreeBSD är intresserad av att få saker gjorda, ochinte emot skada människor som får i deras väg.<Hoponpop> NetBSD är intresserad av att se ingenting blir gjort, och           inte emot skada människor som försöker åstadkomma saker.<Hoponpop> OpenBSD är intresserad av att titta bra, och inte skadar någon           i sin egen lilla samhället, men ser ut alla andra!
		-- David Leimbach

%
<Liiwi> så, vad är det officiella sättet att få buildd att försöka igen ett paket? prod        den med en pinne?<Joey> prod neuro<Liiwi> med en pinne?<Joey> ja.
		-- David Leimbach

%
<Knghtbrd> "... du kommer mer än sannolikt se alla typer av kompilatorn           varningar rulla förbi på skärmen. Detta är normalt och kanvara ignoreras. "<LordHavoc> Knghtbrd: är att en anteckning fäst vid vissa M $ kod?<Knghtbrd> Nej, det är en anteckning om ett gäng GNU saker.
		-- David Leimbach

%
<Hydroxide> knightbrd: från knightbrd.brain import * :)<Knghtbrd> Oh gudar om det vore så enkelt ..<Knghtbrd> från carmack.brain import OpenGL
		-- David Leimbach

%
<LIM> mmmm, multitextured munkar ....<Knghtbrd> LIM: med fruktfyllning?<LIM> knghtbrd: chokladkräm ...
		-- David Leimbach

%
<StevenK> Du skriva delar av Quake i * Python *?<Knghtbrd> MUAHAHAHA
		-- David Leimbach

%
## A_nick (nobody@c213-89-87-111.cm-upc.chello.se) har gått #python<A_nick> Hur lägger jag till en ny nyckel till ett lexikon?<A_nick> nm<Streck> heh :)<Streck> skåda problemlösning makt #python.
		-- David Leimbach

%
<Hop_> jag hade något som jag tror var kyckling som var belagd med en röd       pasta som verkade bestå av lut baseras på hur mycket av min       Tounge det bränns bort.<Hop_> vår vän som är indiska sade att detta är varför de flesta indianer är tunna       och jag citerar "Det tar inte så mycket av denna mat för att få dig       nöjda enoguh att sluta äta. "
		-- David Leimbach

%
<Avsikt> "Det är klassiska sippra upp ekonomi, som erkänner att pengar            är som gödsel: Det fungerar bäst om du sprida det runt ".<Knghtbrd> Avsikt: Carters korrelation: Personer med massor av antingen           vanligen luktar roligt<Avsikt> Knghtbrd: Du SO vinna.
		-- David Leimbach

%
