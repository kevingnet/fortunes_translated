En Linux-maskin! eftersom en 486 är en fruktansvärd sak att avfall!(Genom jjs@wintermute.ucr.edu, Joe Sloan)
		-- Ronald Florence <ron@18james.com> in

%
"Absolut ingenting bör ingås av dessa siffror med undantag av attInga slutsatser kan dras från dem. "(Av Joseph L. Brothers, Linux / PowerPC Project)
		-- Ronald Florence <ron@18james.com> in

%
Egentligen skriva slumpmässiga strängar i Finder gör motsvarandefilnamnskomplettering.(Diskussionen i comp.os.linux.misc på intuition kommandon: filavslutad vs Mac Finder.)
		-- Ronald Florence <ron@18james.com> in

%
Efter att ha sett min nyligen pensionerad pappa tillbringar två veckor att lära sig hur man gör en nymapp, blev det uppenbart att "intuitiv" mestadels betyder "vad författaren ellerhögtalare intuitiva gillar ".(Bruce Ediger, bediger@teal.csn.org i comp.os.linux.misc på xintuition av en Mac-gränssnittet.)
		-- Ronald Florence <ron@18james.com> in

%
"Alla designers språk arrogant. Går med territorium ..."(Av Larry Wall)
		-- Ronald Florence <ron@18james.com> in

%
Och 1.1.81 är officiellt Bugffri (tm), så om du får någon bugg-rapporterpå det, du vet att de är bara onda lögner. "(Av Linus Torvalds, Linus.Torvalds@cs.helsinki.fi)
		-- Ronald Florence <ron@18james.com> in

%
"... Och lättklädda kvinnor, naturligtvis. Vem bryr sig om det är minusgraderutanför"(Av Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
"Och nästa gång du överväga att klaga att köra Lucid Emacs19.05 via NFS från en avlägsen Linux-maskin i Paraguay verkar intefå bakgrundsfärger rätt, vet du vem du ska tacka. "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
>: Alla bärare ute ska känna gladare veta att december är sjöfarten>: Mig en AlphaPC som jag har för avsikt att försöka få Linux körs på: detta kommer>: Definitivt hjälpa spola ut några av de mest flagranta oportabla saker.>: Alpha är mycket mer annorlunda än i386 än 68k saker är, så>: Det är sannolikt att få de flesta av de saker fast.>> Det är inlägg som detta som nästan övertyga oss icke-troende att det> Verkligen är en gud.(En uppföljning av alovell@kerberos.demon.co.uk, Anthony Lovell, till Linusanmärkningar om portering)
		-- Ronald Florence <ron@18james.com> in

%
Den som tror UNIX är intuitiv ska tvingas skriva 5000 raderkod med ingenting men vi eller Emacs. AAAAACK!(Diskussionen i comp.os.linux.misc på intuitiveness kommandon, särskiltEmacs.)
		-- Ronald Florence <ron@18james.com> in

%
"Är [Linux användare] lämlar kollektivt hoppa ut från klippantillförlitlig, väl konstruerad kommersiell programvara? "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
Som vanligt, detta är en 1.3.x release, jag har inte ens sammanställt dennakernel ännu. Så om det fungerar, bör du vara dubbelt imponerad.(Linus Torvalds, meddelar kärnan 1.3.3 på sändlistan linux-kernel.)
		-- Ronald Florence <ron@18james.com> in

%
Undvika helvetets portar. Använd Linux(Okänd källa)
		-- Ronald Florence <ron@18james.com> in

%
Varnas för att skriva \ fBkillall \ fIname \ fP inte kan ha den önskadeeffekt på icke-Linux-system, särskilt när det görs av en privilegierad användare.(Från killall manualsidan)
		-- Ronald Florence <ron@18james.com> in

%
"Dessutom, tror jag [Slackware] låter bättre än" Microsoft ", eller hur?"(Av Patrick Volkerding)
		-- Ronald Florence <ron@18james.com> in

%
Men vad kan man göra med det? - Allestädes närvarande ifrån Linux-användare partner.(Framlagt av Andy Pearce, ajp@hpopd.pwd.hp.com)
		-- Ronald Florence <ron@18james.com> in

%
"Genom golly, jag börjar tro att Linux verkligen * är * det bästa sedanskivat bröd."(Av Vance Petree, Virginia Power)
		-- Ronald Florence <ron@18james.com> in

%
/ * * Oj. Kärnan försökte få tillgång till vissa dåliga sida. Vi måste * Avsluta saker med extrem fördomar.* /die_if_kernel ( "Oj", regs, error_code);(Från linux / arch / i386 / mm / fault.c)
		-- Ronald Florence <ron@18james.com> in

%
"... Djupt Hack Mode - det mystiska och skrämmande tillstånd avmedvetande där Mortal Användare fruktar att beträda. "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
Dijkstra hatar förmodligen mig(Linus Torvalds i kernel / sched.c)
		-- Ronald Florence <ron@18james.com> in

%
DOS: n, en liten irriterande boot virus som orsakar slumpmässigt spontan systemet.     kraschar, oftast bara innan du sparar ett jätteprojekt. Lätt botas genom     UNIX. Se även MS-DOS, IBM-DOS, DR-DOS.(Från David Vickers s .plan)
		-- Ronald Florence <ron@18james.com> in

%
/ * * [...] Observera att 120 sek definieras i protokollet som den maximala * Möjlig RTT. Jag antar att vi måste använda något annat än TCP * Att prata med University of Mars. * TASSAR tillåter oss längre timeout och stora fönster, så när de har genomförts * Ftp till mars kommer att fungera fint. * /(Från /usr/src/linux/net/inet/tcp.c, om RTT [återutsändning timeout])
		-- Ronald Florence <ron@18james.com> in

%
"Ännu mer häpnadsväckande var insikten att Gud har tillgång till Internet. Iundrar om han har en hel nyhetsflöde? "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
> Någonsin hört talas om .cshrc?Det är en stad i Bosnien. Höger?(Diskussionen i comp.os.linux.misc på intuition av kommandon.)
		-- Ronald Florence <ron@18james.com> in

%
Allvarligt fel: Hittade [MS-Windows] System -> Partitionera disk för Linux ...(Genom cbbrown@io.org, Christopher Browne)
		-- Ronald Florence <ron@18james.com> in

%
Hur gör jag skriver "for i in * .dvi gör xdvi jag gjort" i ett GUI?(Diskussionen i comp.os.linux.misc på intuition gränssnitt.)
		-- Ronald Florence <ron@18james.com> in

%
"Hur ska jag veta om det fungerar? Det är vad betatestare är för. Jag barakodad det. "(Skriven Linus Torvalds, någonstans i ett inlägg)
		-- Ronald Florence <ron@18james.com> in

%
---- == - _ / \ /--- == --- (_) __ __ ____ __ / / / \ \- == --- / / _ \ / // / \ \ / / / / _ / \ \ \- ===== / _ / _ // _ / \ _ _ / / _ / \ _ \ / ______ \ \ \En stolt medlem av TeamLinux \ _________ \ /(Genom Chaley (HAC), haley@unm.edu, ch008cth@pi.lanl.gov)
		-- Ronald Florence <ron@18james.com> in

%
Jag utvecklar för Linux för en levande, jag används för att utveckla för DOS.Att gå från DOS till Linux är som handel en segelflygplan för en F117.(Genom entropy@world.std.com, Lawrence Foard)
		-- Ronald Florence <ron@18james.com> in

%
Jag gjorde detta "orsaka Linux ger mig en träig. Det är inte generera intäkter.(Dave '-ddt->' Taylor, meddelar DOOM för Linux)
		-- Ronald Florence <ron@18james.com> in

%
Tveka inte att kontakta mig (flammar om min engelska och värdelös i dennaFöraren kommer att omdirigeras till / dev / null, oh nej, det är fullt ...).(Michael Beck, beskriver PC-högtalare ljudenhet)
		-- Ronald Florence <ron@18james.com> in

%
"Jag vet inte varför, men första C-program tenderar att se en mycket värre änförsta programmen på något annat språk (kanske med undantag för Fortran, men sedanJag misstänker att alla Fortran program ser ut som `firsts") "(Av Olaf Kirch)
		-- Ronald Florence <ron@18james.com> in

%
"Jag en gång bevittnat en långrandig, månadslånga gräl över användningen avmöss kontra trackballs ... Det var mycket dumt. "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
Jag hävdar fortfarande den grad att utforma en monolitisk kärna 1991 är engrundfel. Var tacksam du är inte min elev. Du skulle inte få enhögvärdigt för en sådan konstruktion :-)(Andrew Tanenbaum till Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
"Jag skulle hellre tillbringar 10 timmar att läsa någon annans källkod än10 minuter att lyssna på musak väntar för teknisk support som inte är det. "(Med Dr Greg Wettstein, Roger Maris Cancer Center)
		-- Ronald Florence <ron@18james.com> in

%
"Jag skulle krypa över ett tunnland av" Visual Detta ++ "och" Integrerad utvecklingDet för att komma till gcc, Emacs, och GDB. Tack."(Av Vance Petree, Virginia Power)
		-- Ronald Florence <ron@18james.com> in

%
"Jag är en idiot .. Åtminstone här [bug] tog ca 5 minuter för att hitta .."(Linus Torvalds som svar på en felrapport.)> Jag är en idiot .. Åtminstone [bug] tog ca 5 minuter för att hitta ..Oroande ...(Gonzalo Tornaria som svar på Linus Torvalds: s utskick om en kärna bugg.)> Jag är en idiot .. Åtminstone [bug] tog ca 5 minuter för att hitta ..Vi måste hitta några nya termer för att beskriva resten av oss vanliga dödligasedan.(Craig Schlenter som svar på Linus Torvalds: s utskick om en kärna bugg.)> Jag är en idiot .. Åtminstone [bug] tog ca 5 minuter för att hitta ..Visst, är Linus talar om vilken typ av idioti som andra strävar efter att :-).(Bruce Perens som svar på Linus Torvalds: s utskick om en kärna bugg.)
		-- Ronald Florence <ron@18james.com> in

%
Jag har kört DOOM mer i de senaste dagarna än vad jag har de sistamånader. Jag älskar bara felsökning ;-)(Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
Microsoft Corp., som berörs av den växande populariteten för den fria 32-bitarsoperativsystem för Intel-system, Linux, har anställt ett antal toppprogrammerare från den underjordiska världen av virus utveckling. Bill Gates uppgavigår: "Världsdominans, snabb - det är antingen oss eller Linus". Mr Torvaldsvar inte tillgänglig för en kommentar ...(Rjm@swift.eng.ox.ac.uk (Robert Manners), i comp.os.linux.setup)
		-- Ronald Florence <ron@18james.com> in

%
    if (argc> 1 && strcmp (argv [1], "-Råd") == 0) {printf ( "Do not Panic \ n");exit (42);    }(Arnold Robbins i LJ februari '95, beskriver RCS)
		-- Ronald Florence <ron@18james.com> in

%
+ # Om definitionen (__ alpha__) && definierade (CONFIG_PCI)+ / *+ * Meningen med livet, universum och allting. Plus+ * Detta gör år blir rätt.+ * /+ År - = 42;+ # Endif(Från plåstret för 1.3.2: (kärna / time.c), framlagt av Marcus Meissner)
		-- Ronald Florence <ron@18james.com> in

%
"Om framtida navigationssystem [för interaktiva nättjänster påNII] ser ut som något från Microsoft, kommer det aldrig att fungera. "(Ordförande för Walt Disney Television & telekommunikation)
		-- Ronald Florence <ron@18james.com> in

%
"Om du vill resa runt i världen och bli inbjuden att tala på en hel delolika platser, bara skriva ett Unix-operativsystem. "(Av Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
"[I" Doktor "-läge] Jag tillbringade en bra tio minuter berättar Emacs vad jagtänkte på det. (Svaret var, "Kanske kan du försöka att vara mindremissbruk. ') "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
I de flesta länder som säljer skadliga saker som droger är straffbart.Då howcome människor kan sälja Microsofts program och ostraffat?(Genom hasku@rost.abo.fi, Hasse Skrifvars)
		-- Ronald Florence <ron@18james.com> in

%
Intel teknik verkar ha misheard intel marknadsföringsstrategi. Frasenvar "Dela och erövra" inte "Dela och cock upp"(Genom iialan@www.linux.org.uk, Alan Cox)
		-- Ronald Florence <ron@18james.com> in

%
"Det är Gud. Nej, inte Richard Stallman, eller Linus Torvalds, men Gud."(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
LILO, har du mig på mina knän!(Från David Black, dblack@pilot.njin.net, med ursäkter till Derek ochDomino, och Werner Almsberger)
		-- Ronald Florence <ron@18james.com> in

%
Linux är föråldrad(Andrew Tanenbaum)
		-- Ronald Florence <ron@18james.com> in

%
"Linux utgör en verklig utmaning för dem med smak för senthacka (och / eller samtal med Gud). "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
Linux! Gerilla UNIX Development Venimus, Vidimus, Dolavimus.(Genom mah@ka4ybr.com, Mark A. Horton KA4YBR)
		-- Ronald Florence <ron@18james.com> in

%
"... [Linux] förmåga att prata via något medium utom röksignaler."(Med Dr Greg Wettstein, Roger Maris Cancer Center)
		-- Ronald Florence <ron@18james.com> in

%
linux: därför att en PC är ett ruskigt ting till(Ksh@cis.ufl.edu sätta detta på tshirts i '93)
		-- Ronald Florence <ron@18james.com> in

%
Linux: Eftersom en dator är en fruktansvärd sak att avfall.(Genom komarimf@craft.camp.clarkson.edu, Mark Komarinski)
		-- Ronald Florence <ron@18james.com> in

%
linux: valet av en GNU generation(Ksh@cis.ufl.edu sätta detta på tshirts i '93)
		-- Ronald Florence <ron@18james.com> in

%
"Linux: operativsystemet med en ledtråd ...Command Line användarmiljö ".(Sett i ett inlägg i comp.software.testing)
		-- Ronald Florence <ron@18james.com> in

%
lp1 i brand(En av de mer förvrängd meddelandena från kärnan)
		-- Ronald Florence <ron@18james.com> in

%
Microsoft är inte svaret.Microsoft är frågan.NEJ (eller Linux) är svaret.(Taget från en .signature från någon från Storbritannien, källa okänd)
		-- Ronald Florence <ron@18james.com> in

%
'Mounten' wird fuer drei Dinge benutzt: 'Aufsitzen' auf Pferde, 'einklinken'von Festplatten i Dateisysteme, und, nunna, "besteigen" beim Sex.(Christa Keil i en tysk inlägg: "Montering används för tre saker:klättrar på en häst, som förbinder i en hårddiskenhet i datasystem, och, ja,montering under sex ".)
		-- Ronald Florence <ron@18james.com> in

%
"MSDOS inte få så illa som det är över en natt - det tog över tio årnoggrann utveckling. "(Med dmeggins@aix1.uottawa.ca)
		-- Ronald Florence <ron@18james.com> in

%
"Gör aldrig några mistaeks."(Anonymous, i ett mail diskussion om en kärna felrapport.)
		-- Ronald Florence <ron@18james.com> in

%
Inte jag, killen. Jag läste Bash man sidan varje dag som ett Jehovas vittne läserBibeln. Nej vänta, Bash man page är Bibeln. Ursäkta mig...(Mer om förvirrande alias, tas från comp.os.linux.misc)
		-- Ronald Florence <ron@18james.com> in

%
"Observera att om jag kan få dig att \" SU och säga \ "något bara genom att fråga,du har en mycket allvarlig säkerhets problem på ditt system och du börundersöka saken. "(Av Paul Vixie, vixie-cron 3.0.1 installations anteckningar)
		-- Ronald Florence <ron@18james.com> in

%
Nu vet jag någon där ute kommer att hävda, "Nå, är UNIX intuitiv,eftersom du bara behöver lära 5000 kommandon och sedan allt annat följerfrån det! Har har har! "(Andy Bates i comp.os.linux.misc på "intuitiva", någotförsvara Mac.)
		-- Ronald Florence <ron@18james.com> in

%
Nu är det vi hade den här sortens saker:  ge -a för avkastning till all trafik  ge -t för avkastning på lastbilar  ge -f för avkastning till människor som gick (utbyte fot)  ge -d t * för avkastning på dagar som börjar med t... Du skulle ha en massa döda människor i korsningar och trafikstockningar duskulle inte tro ...(Diskussionen i comp.os.linux.misc på intuition av kommandon.)
		-- Ronald Florence <ron@18james.com> in

%
"På en normal ascii linje, är det enda säkra villkor för att upptäcka en" rast "- Allt annat har tilldelats funktioner genom GNU Emacs ".(Genom Tarl Neustaedter)
		-- Ronald Florence <ron@18james.com> in

%
"På Internet, ingen vet du använder Windows NT"(Framlagt av Ramiro Estrugo, restrugo@fateware.com)
		-- Ronald Florence <ron@18james.com> in

%
En gång i tiden fanns det en DOS användare som såg Unix, och såg att det varbra. Efter att skriva cp på sin DOS maskin hemma, hämtade han GNU sUNIX-verktyg portas till DOS och installerat dem. Han rm'd, cp'd och mv'dLyckligtvis för många dagar, och på att hitta elvis, vi'd han och var glad. Efteren lång dag på jobbet (på en Unix box) han kom hem, började redigera en fil,och kunde inte räkna ut varför han inte kunde avbryta vi (w / ctrl-z) att göraen kompilera.(Genom ewt@tipper.oit.unc.edu (Erik Troan)
		-- Ronald Florence <ron@18james.com> in

%
>> Andra än det faktum Linux har ett coolt namn, kan någon förklara varför jag>> Bör använda Linux över BSD?>> Nej, det är det. Den svala namn, är det. Vi har arbetat mycket hårt på> Skapa ett namn som skulle tilltala de flesta människor, och det> Verkligen lönat sig: tusentals människor använder Linux bara för att kunna> Att säga "OS / 2? Hah. Jag har Linux. En sval namn". 386bsd gjorde> Misstaget att sätta en massa siffror och konstiga förkortningar i> Namn, och skrämma bort en massa människor bara för att det låter för> Tekniskt.(Linus Torvalds "uppföljning av en fråga om Linux)
		-- Ronald Florence <ron@18james.com> in

%
Personligen tror jag att mitt val i mostest-superlativ-dator krig måstevara HP-48-serien av miniräknare. De kommer att köra nästan vad som helst. Och om dekan inte, medan jag bara koppla in en Linux-burk till den seriella porten och ladda uppHP-48 VT-100 emulatorn.(Genom jdege@winternet.com, Jeff Dege)
		-- Ronald Florence <ron@18james.com> in

%
Det finns inga trådar i a.b.p.erotica, så det finns ingen vinst i att använda engängade nyhetsläsare.(Okänd källa)
		-- Ronald Florence <ron@18james.com> in

%
"Problemlösning under Linux har aldrig varit cirkusen att det är underAIX. "(Av Pete Ehlke i comp.unix.aix)
		-- Ronald Florence <ron@18james.com> in

%
avslutas när sluta uttalande läsa, BC-processor       avslutas, oavsett var avsluta uttalande       ning hittas. Till exempel, "if (0 == 1) quit"       kommer att orsaka bc att avsluta.(Sett på manualsidan för "bc". Notera den "om" uttalande logik)
		-- Ronald Florence <ron@18james.com> in

%
Windows på en Pentium är som att ha en helt ny Porsche men barakunna köra bakåt med handbromsen på.(Okänd källa)
		-- Ronald Florence <ron@18james.com> in

%
"Sic transit discus mundi"(Från systemadministratörer, av Lars Wirzenius)
		-- Ronald Florence <ron@18james.com> in

%
Suck. Jag vill gärna tro att det är bara Linux människor som vill vara påden "framkant" så illa att de går direkt från stupet.(Craig E. Groeschel)
		-- Ronald Florence <ron@18james.com> in

%
Den chattprogram är i offentligt område. Detta är inte den offentliga licensen GNU. OmDet bryter då du får behålla båda delar.(Upphovsrätts för chattprogram)
		-- Ronald Florence <ron@18james.com> in

%
> Dagen människor tror Linux skulle vara bättre betjänt av någon annan (FSF> Är det naturliga alternativet), jag kommer "abdikera". Jag tror inte att> Det är något folk har att oroa sig för just nu - Jag ser inte det> Händer inom en snar framtid. Jag gillar att göra Linux, även om det gör> Innebär en del arbete, och jag har inte fått några klagomål (vissa nästan skygg> påminnelser om en lapp jag har glömt eller ignoreras, men ingenting> Negativt hittills).>> Ta inte ovan att innebära att jag ska sluta dagen någon klagar:> Jag är okänslighet (Lasu, som läser detta över min axel kommenterade> Som "tjock-headed är närmare sanningen") nog att ta lite missbruk.> Om jag inte var, skulle jag har slutat att utveckla Linux dagen ast förlöjligade mig> Om c.o.minix. Vad jag menar är bara att medan Linux har mitt barn så> Långt, jag vill inte stå i vägen om man vill göra något> Bättre av det (*).>> Linus>> (*) Hej, jag kanske skulle kunna ansöka om ett helgon-hood från påven. gör> Någon vet vad hans e-postadress är? Jag är så trevligt det gör du puke.(Utdrag ur Linus svar på någon orolig för framtiden för Linux)
		-- Ronald Florence <ron@18james.com> in

%
Det fina med Windows är - Det är inte bara kraschar, det visar endialogrutan och låter du trycker på "OK" först.(Arno Schaefer s .sig)
		-- Ronald Florence <ron@18james.com> in

%
Den enda "intuitiva" gränssnitt är bröstvårtan. Efter det är det alla lärt.(Bruce Ediger, bediger@teal.csn.org i comp.os.linux.misc på X-gränssnitt.)
		-- Ronald Florence <ron@18james.com> in

%
Det finns två typer av Linux-utvecklare - de som kan stava, ochde som inte kan. Det finns en konstant fältslag mellan de två.(Från en av de efter 1.1.54 kärna uppdateringsmeddelanden skickas till c.o.l.a)
		-- Ronald Florence <ron@18james.com> in

%
Det här meddelandet skickades av Linux, den fria Unix.Windows utan X är som att älska utan en partner.Sex, Drugs & Linux reglerwin-nt från de människor som uppfann Edlinäpplen har inneburit problem sedan edenLinux, sättet att bli av med boot virus(Genom mwikholm@at8.abo.fi, Madsen Wikholm)
		-- Ronald Florence <ron@18james.com> in

%
"... Unix, MS-DOS och Windows NT (även känd som den gode, den onde, ochden fula)."(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
"... Mycket få fenomen kan dra någon ur djup Hack läge med tvånoterade undantag: att träffas av blixten, eller ännu värre, din * dator *att träffas av blixten. "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
"Vinka bort ett moln av rök, jag ser upp, och är förblindade av en ljus, vitljus. Det är Gud. Nej, inte Richard Stallman, eller Linus Torvalds, men Gud. Ien blomstrande röst, säger han: "Detta är ett tecken använder Linux, den fria UNIX-system.FÖR 386. "(Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
"Vi vet alla Linux är stor ... det gör oändliga loopar i 5 sekunder."(Linus Torvalds om överlägsenheten av Linux på AmsterdamLinux Symposium)
		-- Ronald Florence <ron@18james.com> in

%
Vi är Microsoft. Du kommer att assimileras. Motstånd är meningslöst.(Skriven B.G., Gill Bates)
		-- Ronald Florence <ron@18james.com> in

%
Vi är Pentium Borg. Division är meningslöst. Du kommer att approximeras.(Sett i någons .signature)
		-- Ronald Florence <ron@18james.com> in

%
Vi använder Linux dagligen till UPP produktiviteten - så upp din!(Anpassad från Pat Paulsen av Joe Sloan)
		-- Ronald Florence <ron@18james.com> in

%
Vi kommer att begrava DOS, inte att berömma det.(Paul Vojta, vojta@math.berkeley.edu, omskriva ett citat av Shakespeare)
		-- Ronald Florence <ron@18james.com> in

%
Vi använder Linux för alla våra verksamhetskritiska applikationer. Med källkodeninnebär att vi inte hålls som gisslan av någon supportavdelning.(Russell Nelson, VD för Crynwr Software)
		-- Ronald Florence <ron@18james.com> in

%
"Vad du sluta med, efter att ha kört ett operativsystem koncept genommånga marknadsföring kaffefilter, är något som inte till skillnad från vanlig varmvatten."(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
Vad detta script göra?    packa upp; Rör ; finger; mount; gasp; ja; umount; sovaTips för svaret: inte allt är datororienterade. Ibland är dui en sovsäck, camping.(Bidrag från Frans van der Zande.)
		-- Ronald Florence <ron@18james.com> in

%
'När du säger "Jag skrev ett program som kraschat Windows", människor bara stirrar pådu uttryckslöst och säga "Hej, jag fick de med systemet, * gratis *". "(Av Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
"Piska mig. Slå mig. Gör mig upprätthålla AIX."(Av Stephan Zielinski)
		-- Ronald Florence <ron@18james.com> in

%
"Vem är General Failure och varför han läser min hårddisk?"Microsoft spel chekar vor segel, worgs galler !!(Genom leitner@inf.fu-berlin.de, Felix von Leitner)
		-- Ronald Florence <ron@18james.com> in

%
Vem vill komma ihåg att fly-x-alt-kontroll vänster shift-b sätter dig insuper-edit-debug-kompilera läge?(Diskussionen i comp.os.linux.misc på intuitiveness kommandon, särskiltEmacs.)
		-- Ronald Florence <ron@18james.com> in

%
Varför använder Windows, eftersom det finns en dörr?(Genom fachat@galileo.rhein-neckar.de, Andre Fachat)
		-- Ronald Florence <ron@18james.com> in

%
"Världsdominans. Snabb"(Av Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
..du kunde tillbringa * hela dagen * anpassa namnlisten. Tro mig. jagtalar av erfarenhet. "(Av Matt Welsh)
		-- Ronald Florence <ron@18james.com> in

%
"... Kan man lika gärna hoppa över Xmas firandet helt och i ställetsitta framför din Linux-dator spelar medall-new-och-förbättrad Linux-kärnan version. "(Av Linus Torvalds)
		-- Ronald Florence <ron@18james.com> in

%
Ditt jobb är att vara en professor och forskare: Det är ett helvete av en bra ursäktför vissa av de hjärn skador av minix.(Linus Torvalds till Andrew Tanenbaum)
		-- Ronald Florence <ron@18james.com> in

%
Jag har hört en Judisk och en muslim argumentera i en Damaskus café med mindre lidelseän Emacs krig. "<Ueu1c4mbrc.fsf@auda.18james.com>
		-- Ronald Florence <ron@18james.com> in

%
