1/2 oz. gin1/2 oz. vodka1/2 oz. rom (företrädesvis mörk)3/4 oz. tequilla1/2 oz. triple sec1/2 oz. apelsinjuice3/4 oz. sour mix1/2 oz. colaskaka med is och sila upp i frostat glas.Long Island Iced Tea
		-- Dean Martin

%
6 oz. apelsinjuice1 oz. vodka1/2 oz. gallianoHarvey Wallbanger
		-- Dean Martin

%
En öl försenad är en öl förnekas.
		-- Dean Martin

%
Ett par fler skott av whisky, kvinno runt här börjar ser bra ut.[Något om en 10 är en 4 efter en sex-pack? Ed.]
		-- Dean Martin

%
En kille går in i en bar, beställer en öl, bär den på toaletten och dumpar deti en pissoar. Under de närmaste timmarna, går han tillbaka till barenoch upprepar denna sekvens - flera gånger. Slutligen bartendern fick såmärkligt att han lutade sig över baren och frågade honom vad han gjorde.Svarade kunden "Undvika mellanhand."
		-- Dean Martin

%
En förbuds är den sortens människa man inte bryr sig att dricka med- Även om han drack.
		-- H. L. Mencken

%
Absinthe gör tårta växa Fonder.
		-- H. L. Mencken

%
Alkohol är anestesi genom vilken vi uthärda driften av livet.
		-- George Bernard Shaw

%
Alkohol, hasch, blåsyra, stryknin är svaga utspädningar. det säkrastegift är dags.
		-- Emerson, "Society and Solitude"

%
Anonyma Alkoholister är när man får dricka under någon annans namn.
		-- Emerson, "Society and Solitude"

%
Förvara alltid öl på en mörk plats.
		-- Lazarus Long

%
En alkoholist är någon du inte gillar som dricker så mycket som du gör.
		-- Dylan Thomas

%
Och du kan inte få någon Watney Red Barrel,eftersom staplarna stänger varje gång du är törstig ...
		-- Dylan Thomas

%
... Åtminstone jag trodde jag dansade, 'til någon klev på min hand.
		-- J. B. White

%
Var försiktig med starka drycker. Det kan göra dig skjuta på tullindrivare och miss.
		-- Lazarus Long, "Time Enough for Love"

%
Eftersom vinet kommer ihåg.
		-- Lazarus Long, "Time Enough for Love"

%
Öl & kringlor - Frukost of Champions.
		-- Lazarus Long, "Time Enough for Love"

%
Öl - det är inte precis för frukost anymore.
		-- Lazarus Long, "Time Enough for Love"

%
Tiggare till välklädda affärsman:"Kan du avvara $ 20,95 för en femtedel av Chivas?"
		-- Lazarus Long, "Time Enough for Love"

%
Bästa Öl: En panel av provsmakare monteras av konsumentens unionen 1969bedömas Coors och Miller High Life att vara bland de allra bästa. De somtvekan om att öl är ett allvarligt ämne kan begrunda dess effekt på amerikanskahistoria. Till exempel beslutade New Englands första kolonister att ankrapå Plymouth Rock stället för att fortsätta vidare till Virginia eftersom, som en avdem uttryckte det, "Vi kunde inte nu ta tid för vidare behandling, vårproviant spenderas och särskilt vår öl. "
		-- Felton & Fowler's Best, Worst & Most Unusual

%
Sprit är svaret. Jag minns inte frågan.
		-- Felton & Fowler's Best, Worst & Most Unusual

%
bytet konjak-och-vatten två bra saker.
		-- Charles Lamb

%
Men, officer, han är inte druckit, jag såg bara hans fingrar rycka!
		-- Charles Lamb

%
Cerebus: Jag skulle älska att slicka aprikos brandy ur naveln.Jaka: Titta, har Cerebus-- Jaka att berätta ... någotCerebus: Om Cerebus hade en navel, skulle du slicka aprikos brandy ut av det?Jaka: Ugh!Cerebus: Du tycker inte om aprikos brandy?
		-- Cerebus #6, "The Secret"

%
Rödvin är sprit för pojkar; port för män; men han som strävar efter att vara en hjälte... Måste dricka konjak.
		-- Samuel Johnson

%
Klättra upp en barstol, ett snöre bad om en öl."Vänta en minut. Är du en sträng?""Ja, ja, jag är.""Tyvärr. Vi serverar inte strängar här."Den bestämda strängen lämnade baren och stoppade en förbipasserande. "Ursäkt,mig ", det sade," skulle du strimla mina ändar och binda upp mig som en kringla? "Theförbipasserande skyldig, och strängen åter in i baren. "Kan jag få en öl,vänligen? "Det frågade bartendern.Barkeep in en öl framför strängen, sedan plötsligt stannade."Hej, är du inte strängen jag bara kastade ut härifrån?""Nej, jag är en sliten knut."
		-- Samuel Johnson

%
Coach: Kan jag dra dig en öl, Norm?Norm: Nej, jag vet hur de ser ut. Häll mig bara en.Coach: Vad sägs om en öl, Norm?Norm: Hej Jag är hög på livet, tränare. Naturligtvis är öl mitt liv.Coach: Hur är en öl ljud, Norm?Norm: Jag vet inte. Jag brukar avsluta dem innan de får ett ord i.
		-- Cheers, Fortune and Men's Weights

%
Coach: Hur går det, Norm?Norm: Pappa rika och Mommas bra lookin '.Sam: Vad är upp, Norm?Norm: Mina bröstvårtor. Det är kallt ute.Coach: Vad är historien, Norm?Norm: Törstig killen går in i en bar. Du avsluta det.
		-- Cheers, Endless Slumper

%
Tränare: Vad skulle du säga till en öl, Normie?Norm: pappa wuvs dig.Sam: Vad du vill, Normie?Norm: En anledning att leva. Gimme en annan öl.Sam: Vad kommer du att ha, Norm?Norm: Tja, jag är i ett spel humör, Sammy. Jag tar ett glas vad      kommer ut ur den kranen.Sam: Åh, ser ut som öl, Norm.Norm: Kalla mig Mister Lucky.
		-- Cheers, The Executive's Executioner

%
Coach: Vad är upp, Norm?Norm: mungiporna, Coach.Coach: Vad skakar, Norm?Norm: Alla fyra kinder och ett par hakor, tränare.Coach: Öl, Normie?Norm: Öh, tränare, jag vet inte, jag hade en i veckan. Eh, varför inte, jag är fortfarande ung.
		-- Cheers, Snow Job

%
Kom snabbt, jag smaka stjärnor!
		-- Dom Perignon, upon discovering champagne.

%
Kom, hyresvärd, fylla den strömmande skål tills det löper över,Ikväll kommer vi alla glatt vara - i morgon kommer vi att få nykter.
		-- John Fletcher, "The Bloody Brother", II, 2

%
Drick inte när du kör - du kanske slå ett gupp och spilla den.
		-- John Fletcher, "The Bloody Brother", II, 2

%
Rök inte nästa cigarett. Upprepa.
		-- John Fletcher, "The Bloody Brother", II, 2

%
Dryck Canada Dry! Du kanske inte lyckas, men det * __ är * kul att försöka.
		-- John Fletcher, "The Bloody Brother", II, 2

%
Dricka kaffe för omedelbar avkoppling? Det är som att dricka alkohol föromedelbara motorik.
		-- Marc Price

%
Dricka är inte en publiksport.
		-- Jim Brosnan

%
Dricka gör sådana dårar människor, och människor är sådana idioter att börjamed att det förvärrar ett brott.
		-- Robert Benchley

%
Drunks är sällan underhållande om de inte vet några bra låtar och förlorarmycket poker.
		-- Karyl Roosevelt

%
Eggnog är en traditionell semester drink uppfanns av den engelska. Mångafolk undrar där ordet "äggtoddy" kommer från. Den första stavelsenkommer från det engelska ordet "ägg", som betyder "ägg". Jag vet inte varden "nog" kommer ifrån.För att göra äggtoddy, måste du rom, whisky, vin gin och, om de är isäsong, ägg ...
		-- Karyl Roosevelt

%
ELECTRIC JELL-O2 lådor JELL-O varumärke gelatin 2 paket Knox varumärke unflavored gelatin2 koppar frukt (en sort) 2+ dl vatten1/2 flaska Everclear varumärke spritMix JELL-O och Knox gelatin i 2 koppar kokande vatten. Rör 'tilfullständigt upplöst.Häll varma blandningen i en platt panna. (JELL-O formar kommer inte att fungera.)Rör i sprit i stället för vanligt kallt vatten. Ta bort eventuella stelGlops av slem. (Alkohol har en ovanlig effekt på överskott JELL-O.)Häll i frukt till önskad smak, och för att absorbera överskott av alkohol.Blanda i lite kallt vatten för att späda ut alkohol och göra det lättare att äta försvag i hjärtat.Kylskåp över natten för att tillåta blandningen att fullständigt härda. (ca 8-12 timmar.)Skär i rutor och mycket nöje!VARNING:Håll ingredienser borta från öppen eld. rekommenderas inte förbarn under åtta års ålder.
		-- Karyl Roosevelt

%
Varje morgon är en Smirnoff morgon.
		-- Karyl Roosevelt

%
Utmärkt dag för att dricka tungt. Spike kontoret vattenkylare.
		-- Karyl Roosevelt

%
Festnivå 1: Dina gäster chattar vänligt med varandraandra, beundrar dina julgransprydnader, sjunger julsånger runtpianot, smuttar på sina drinkar och knaprar smårätter.Festnivå 2: Dina gäster pratar högljutt - iblandtill varandra, och ibland ingen alls, ordna dinJulgransprydnader, sjunger "I Gotta Be Me" runt upprättpiano, svälja sina drycker och vräker ner smårätter.Festnivå 3: Dina gäster argumenterar våldsamt medlivlösa föremål, sjunger "jag kan inte få någon tillfredsställelse," svälja nerandras drycker, vräker i sig julgransprydnader ochplacera smårätter i piano för att se vad som händer närde små hammare slår.Festnivå 4: Dina gäster, smårätter smort heladeras nakna kroppar utför en rituell dans runt den brinnandeJulgran. Pianot saknas.Du vill behålla din fest någonstans runt nivå 3, såvida intedu hyr din bostad och egna skjutvapen, i vilket fall du kan gå till nivå4. Det bästa sättet att komma till nivå 3 är ägg-nog.
		-- Karyl Roosevelt

%
Fiske, med mig, har alltid varit en ursäkt för att dricka på dagtid.
		-- Jimmy Cannon

%
Fortune avslutar de stora citat, # 17"Denna knopp av kärlek, av sommarens mognad andedräkt,Kan visa sig vara en sköna blomma när nästa vi träffas. "Juliet, är det här knopp för dig.
		-- Jimmy Cannon

%
Fortunes favoritrecept: # 8Christmas Rum Cake1 eller 2 liter rom 1 msk. bakpulver1 kopp smör 1 tsk. soda1 tsk. socker 1 msk. citronjuice2 stora ägg 2 dl farinsocker2 koppar torkad diverse frukt 3 koppar hackade engelska valnötterInnan du börjar prova rom för att kontrollera kvaliteten. Bra, är inte det? NuVälj en stor bunke, mätglaset, etc. Kontrollera rom igen. Detmåste vara precis rätt. Var noga med rom är av högsta kvalitet. Häll en kopprom i ett glas och dricker det så fort som möjligt. Upprepa. Med en elektriskmixer, slå en kopp smör i en stor fluffig skål. Lägga en seaspoon av tugaroch slå igen. Samtidigt se till rom coh absolut högsta kvalitet.Prov en annan kopp. Öppna andra kvart efter behov. Tillsätt 2 orge laggs, 2 kopparstekt druit och slå tills hög. Om stekt druit fastnar ivispar, bara bända loss den med en skruvmejsel. Prov rom igen, kontrollför toncisticity. Nästa sålla 3 koppar bakpulver, en nypa rom, enseaspoon av toda och en kopp peppar eller salt (det egentligen ingen roll).Prova några mer. Sålla 912 pint citronsaft. Vik in schopped smör ochansträngda chups. Lägg bablespoon brun gugar, eller vad färg du har.Blanda mell. Fett ugn och vrid kakform till 350 gredees och rake tillspoothtick kommer ut crean.
		-- Jimmy Cannon

%
FORTUNE parti TIPS # 14Trött på att finna att andra människor att hjälpa sig själva till godasprit vid BYOB partierna? Ta med en ljus, som du sätter ochljus efter att du har öppnat flaskan. Ingen har någonsin förväntar sig någotdrickbart för att vara i en flaska som har ett ljus fastnat i dess hals.
		-- Jimmy Cannon

%
Glögg (en traditionell skandinavisk semester dryck):femtedel av torrt rött vinfemtedel av Aquavit1 och 1/2 tums bit av kanel10 kardemumma frön1 kopp russin4 torkade fikon1 kopp skål eller mandelspånnågra bitar av torkad apelsinskal5 kryddnejlika1/2 lb. sockerbitarVärma upp vin och hårda saker (som kan vara substituerad med vinför svag i hjärtat) i en stor pott efter att ha lagt alla andra saker UTOMsockerbitar. Just när det når kokpunkten, sätta sockret i en trådsil, fukta den i den heta brygd, lyft ut och tända den med en tändsticka.Doppa sockret flera gånger i vätskan tills allt är upplöst. Tjänahet i koppar med några russin och mandel i varje kopp.OBS. Akvavit kan vara svårt att hitta och dyrt för start. Använd det baraom du verkligen har en djupt rotad önskan att vara noga, eller om du är i svenskaextraktion.
		-- Jimmy Cannon

%
Halleys komet: Det kom, vi såg, vi drack.
		-- Jimmy Cannon

%
Harrys bar har en ny cocktail. Det kallas MRS punch. De gör det medmjölk, rom och socker och det är fantastiskt. Mjölken är för vitalitet ochsocker är för pep. De satte i rom så att folk vet vad de ska göramed allt vad det pep och vitalitet.
		-- Jimmy Cannon

%
Att ha en underbar vin, önskar att du var öl.
		-- Jimmy Cannon

%
Efter att ha vandrat löst in i en bländande snöstorm Sam var kraftigtlättad över att se en kraftig St Bernard hund avgränsar mot honom medden traditionella fatet konjak fastspänd på hans krage."Äntligen" ropade Sam "människans bästa vän - och en stor stor hund, också!"
		-- Jimmy Cannon

%
Han kände tavernes väl i varje toun.
		-- Geoffrey Chaucer

%
Han är precis som Capistrano, alltid redo för några klunkar.
		-- Geoffrey Chaucer

%
"Hej! Vem tog korken av min lunch ??!"
		-- W. C. Fields

%
Hogans hjältar dricka spel -Ta ett skott varje gång:- Sergeant Schultz säger: "Jag knoooooowww nooooothing!"- General Burkhalter eller Major Hochstetter skrämma / förolämpning överste Klink.- Överste Klink faller för överste Hogan smicker.- En av fångarna smyger ut ur lägret (ett skott för varje fånge att gå).- Överste Klink snaps till uppmärksamhet efter att svara i telefon (två skottom det är en av våra hjältar i den andra änden).- En av tyskarna hotas med att skickas till den ryska fronten.- Korpral Newkirk kallar upp en tysk i sin bluff tysk accent, ochtricks honom (två skott om det är överste Klink).- Hogan har en romantisk mellanspel med en vacker flicka från tunnelbanan.- Överste Klink berättar hur han aldrig har haft en flykt från Stalag 13.- Sergeant Schultz ger upp en hemlig (två skott om han mutade med mat).- Fångarna lyssna på tyskarnas samtal med en dold sändare.- Sergeant Schultz "fångar" en av fångarna efter en flykt.- Lebeau uttalar "överste" som "CUH-loh-`nell".- Carter bygger någon form av anordning (två skott om det inte är explosivt).- Lebeau bär hans förkläde.- Hogan säger: "Vi har inget annat val" när någon hävdar att planen äromöjligt.
		-- The prisoners capture an important German, and sneak him out the tunnel.

%
Jag kan inte dö förrän regeringen finner en säker plats att begrava min lever.
		-- Phil Harris

%
Jag misstror en man som säger när. Om han måste vara noga med att inte drickaalltför mycket, beror det på att han inte är att lita på när han gör.
		-- Sidney Greenstreet, "The Maltese Falcon"

%
Jag dricker inte, jag tycker inte om det, gör det mig att känna alltför bra.
		-- K. Coates

%
Jag dricker för att göra andra människor intressant.
		-- George Jean Nathan

%
Jag gav upp rökning, alkohol och sex. Det var den mest * __________ skrämmande * 20minuter i mitt liv!
		-- George Jean Nathan

%
Jag har bara haft arton whisky i en rad. Jag tror det är ett rekord.
		-- Dylan Thomas, his last words

%
Jag måste tänka svårt att nämna en intressant man som inte dricker.
		-- Richard Burton

%
Jag kysste min första tjej och rökte min första cigarett på samma dag.Jag har inte haft tid för tobak sedan.
		-- Arturo Toscanini

%
Jag kanske inte kan gå, men jag kör från sittande ställning.
		-- Arturo Toscanini

%
Jag måste få ut av dessa våta kläder och in i en torr Martini.
		-- Alexander Woolcott

%
Jag har aldrig sagt alla demokrater var saloonkeepers; vad jag sa var allasaloonkeepers var demokrater.
		-- Alexander Woolcott

%
Jag tar aldrig jobbet hem med mig; Jag lämnar alltid det i vissa bar längs vägen.
		-- Alexander Woolcott

%
Jag antar att om några timmar kommer jag att nyktra till. Det är en sådan sorgligtyckte. Jag tror att jag kommer att ha några fler drinkar att förbereda mig.
		-- Alexander Woolcott

%
Jag brukade ha en alkoholproblem. Nu älskar jag saker.
		-- Alexander Woolcott

%
Jag kommer inte att dricka!Men om jag gör ...Jag kommer inte att bli full!Men om jag gör ...Jag kommer inte offentligt!Men om jag gör ...Jag kommer inte att falla ner!Men om jag gör ...Jag kommer att falla framsidan nedåt så att de inte kan se mitt företag emblem.
		-- Alexander Woolcott

%
Jag önskar att du var en Scotch on the rocks.
		-- Alexander Woolcott

%
Jag skulle vilja träffa killen som uppfann öl och se vad han arbetar på nu.
		-- Alexander Woolcott

%
Jag vill hellre ha en gratis flaska framför mig än en prefrontala lobotomi.[Också tillskrivas S. Clay Wilson. Ed.]
		-- Fred Allen

%
Jag är inte under alkafluence av inkaholatt vissa thinkle peep jag.Det är bara fullare jag sitta här längre får jag.
		-- Fred Allen

%
Jag har alltid tyckte synd om människor som inte dricker - kom ihåg,när de vaknar, det är så bra som de är gonna känner hela dagen!
		-- Fred Allen

%
Jag har alltid gjort det en högtidlig praxis att aldrig dricka något starkareän tequila innan frukost.
		-- R. Nesson

%
Jag har aldrig varit berusade, men ofta jag har overserved.
		-- George Gobel

%
Om Gud hade tänkt Man Smoke, skulle han ha satt honom på Fire.
		-- George Gobel

%
Om Gud hade tänkt Män Smoke, skulle han ha lagt skorstenar i deras huvuden.
		-- George Gobel

%
Om jag visste vad varumärket [whisky] han dricker, skulle jag skicka ett fat ellerså att mina andra generaler.
		-- Abraham Lincoln, on General Grant

%
Om folk drack bläck i stället för Schlitz, skulle de vara bättre.[Vilket märke av bläck? Ed.]
		-- Edward E. Hippensteel

%
Om du inte dricker det, någon annan kommer.
		-- Edward E. Hippensteel

%
Om du dricker, inte parkera. Olyckor gör människor.
		-- Edward E. Hippensteel

%
År 1967, den sovjetiska regeringen präglat en vacker silver rubel med Lenini en mycket bekant pose - armar ovanför honom, leder landetrotation. Men det var klart för alla, att om du tittat på det frånbakom, var det tydligt att Lenin pekade på 11:00, när vodkabutiker öppnas, och var faktiskt säger, "Kamrater, fram till Vodka butiker.Det blev på modet, när man ville ha en drink, att ta utrubel och säger: "Åh herregud, kamrater, säger Lenin mig att vi bör gå.
		-- Edward E. Hippensteel

%
I en flaska, är halsen alltid överst.
		-- Edward E. Hippensteel

%
I en samling av två eller flera personer, när en tänd cigarett ärplaceras i en askkopp, kommer röken waft in i ansiktet på den icke-rökare.
		-- Edward E. Hippensteel

%
I en whisky det är ålder, i en cigarett det smak och i en sportbildet är omöjligt.
		-- Edward E. Hippensteel

%
I vino veritas.[I vin finns det sanning.]
		-- Pliny

%
Det har sagts att PR är konsten att vinna vänneroch få människor under påverkan.
		-- Jeremy Tunstall

%
Det är en modig man som när det är som mörkast, kan luta sig tillbaka och party!
		-- Dennis Quaid, "Inner Space"

%
Det kommer att bli bra,Det är nästan midnatt,Och jag har två flaskor vin.
		-- Dennis Quaid, "Inner Space"

%
Det är samma gamla historia; pojke möter öl, dricker pojke öl ... pojke fåren annan öl.
		-- Cheers

%
Det är meningslöst att försöka hålla vissa människor att allt de säger när de ärkär i, berusade, eller köra för kontor.
		-- Cheers

%
Håll Amerika vacker. Svälj ölburkar.
		-- Cheers

%
Kiss en icke-rökare, smaka skillnaden.
		-- Cheers

%
Kyssa en rökare är som att slicka en askkopp.
		-- Cheers

%
Lady Astor gav en kostym boll och Winston Churchill frågade henne vadförklädnad hon skulle rekommendera för honom. Hon svarade: "Varför kommer du intenykter, Mr. statsminister? "
		-- Cheers

%
Låt värdiga medborgare Chicago få sin sprit på bästa sättDom kan. Jag är trött på jobbet. Det är en otacksam en och full av sorg.
		-- Al Capone

%
Livet, som öl, är bara lånat.
		-- Don Reed

%
Titta på det här sättet: Din dotter just heter färskt kalkon du toghem "Omfamningar", så att du går ut för att köpa en burk skinka. Och du är fortfarandedricka vanlig scotch?
		-- Don Reed

%
Titta på det här sättet: Din fru spendera 280 $ i månaden på meditation lärdglömma $ 26.000 av högskoleutbildning. Och du fortfarande dricker vanlig scotch?
		-- Don Reed

%
Marvin den naturspionerade en gräshoppa hoppande tillsammans i gräset,och på humör för med naturen, sällsynta även bland fullfjädradNaturälskare, talade han till gräshoppa, säger: "Hej, vängräshoppa. Visste du att de har namngett en drink efter dig? ""Verkligen?" svarade gräshoppa, uppenbarligen nöjd. "De harnamngav en drink Fred? "
		-- Don Reed

%
"Sinne om jag röker?""Jag bryr mig inte om du fattade eld och dö!"
		-- Don Reed

%
"Sinne om jag röker?""Ja, jag skulle vilja se att, det kommer ut ur öronen eller vad?"
		-- Don Reed

%
Min mamma dricker för att glömma hon dricker.
		-- Crazy Jimmy

%
Min morbror var staden full - och vi bodde i Chicago.
		-- George Gobel

%
försena aldrig slutet på ett möte eller början på en cocktail timme.
		-- George Gobel

%
dricker aldrig från fingret skål - det innehåller bara vatten.
		-- George Gobel

%
Nej, jag har inte ett alkoholproblem.Jag dricker, jag bli full, jag faller ner.Inga problem!
		-- George Gobel

%
[Norm kommer in med en attraktiv kvinna.]Coach: Normie, Normie, kan detta vara Vera?Norm: Med en massa dyr operation, kanske.Coach: Vad är upp, Normie?Norm: Temperaturen under min krage, Coach.Tränare: Vad skulle du säga till en trevlig öl, Normie?Norm: Going down?
		-- Cheers, Diane Meets Mom

%
[Norm går in i baren på Vic Bowl-A-Rama.]Utanför skärmen publiken: normen!Sam: Hur fan vet de honom här?Cliff: Han har fått ett liv, du vet.Woody: Vad kan jag göra för dig, mr Peterson?Norm: rymma med min fru.Woody: Hur liv, mr Peterson?Norm: Åh, jag väntar på filmen.
		-- Cheers, Take My Shirt... Please?

%
[Norm är arg.]Woody: Vad vill du ha, mr Peterson?Norm: Clifford Calvin huvud.Sam: Hej, vad som händer, Norm?Norm: Tja, det är en hund-äta-hundvärlden, Sammy,      och jag bär Milk-Bone underkläder.Sam: Hur liv i omkörningsfilen, Normie?Norm: Slår mig, jag kan inte hitta den på rampen.
		-- Cheers, Diane Chambers Day

%
[Norm återvänder från sjukhuset.]Coach: Vad är upp, Norm?Norm: Allt som är tänkt att vara.Sam: Vad är nytt, Normie?Norm: Terrorister, Sam. De har tagit över magen. De kräver öl.Coach: Vad ska det vara, Normie?Norm: Bara vanligt, tränare. Jag har ett skum av öl och en snorkel.
		-- Cheers, King of the Hill

%
[Norm försöker bevisa att han inte är Anton Kreitzer.]Norm: Eftermiddag, alla!All: Anton!Woody: Vad som händer, mr Peterson?Norm: En blinkande skylt i magen som säger, '' Sätt öl här ''.Sam: Vad vill du ha, Norm?Norm: [skrapa skägget] Har någon loppa pulver? Ah, bara skojar.      Gimme en öl; Jag tror att jag bara dränka små rotskott.
		-- Cheers, Two Girls for Every Boyd

%
Norm: Herrar, starta din kranar.Coach: Hur är livet behandlar dig, Norm?Norm: Som det fångade mig i sängen med sin fru.Coach: Hur liv, Norm?Norm: Inte för blödiga, tränare.
		-- Cheers, Friends, Romans, and Accountants

%
Norm: Hej, alla.All: [tystnad; alla är arg på Norm för att vara rik.]Norm: [bär på båda sidor av konversationen själv.]       Norm! (Normand.)       Hur mår du idag, Norm?       Rik och törstig. Häll mig en öl.Woody: Vad är det senaste, mr Peterson?Norm: Zsa-Zsa gifter sig med en miljonär, Peterson dricker en öl.       Film på elva.Woody: Hur mår du idag, Mr. Peterson?Norm: Aldrig varit bättre, Woody. ... Bara en gång skulle jag vilja vara bättre.
		-- Cheers, Chambers vs. Malone

%
Inte alla män som dricker är poeter. Några av oss dricker eftersom vi inte poeter.
		-- Cheers, Chambers vs. Malone

%
Inte dricka, jaga kvinnor, eller göra droger kommer inte att du lever längre -Det verkar bara så.
		-- Cheers, Chambers vs. Malone

%
LÄGGA MÄRKE TILL:Någon sett röka kommer att antas vara i brand och viljasummariskt släcka.
		-- Cheers, Chambers vs. Malone

%
Nu är det dags för att dricka; nu är det dags att slå jorden medohämmad fot.
		-- Quintus Horatius Flaccus (Horace)

%
Naturligtvis elverktyg och alkohol inte blanda. Alla vet maktverktyg är inte lösliga i alkohol ...
		-- Crazy Nigel

%
Gamla farfar är död men hans sprit leva på.
		-- Crazy Nigel

%
När ... i ödemarken i Afghanistan, förlorade jag min korkskruv, och vi vartvingas leva på något annat än mat och vatten i flera dagar.
		-- W. C. Fields, "My Little Chickadee"

%
En skillnad mellan en man och en maskin är att en maskin är tystnär väl oljad.
		-- W. C. Fields, "My Little Chickadee"

%
En dammig juli eftermiddag, någonstans kring sekelskiftet, PatrickMalone var i Mulcahey s Bar, böja en armbåge med den andra gatan bilenledare från Brooklyn Traction Company. Medan de diskuteradefördelarna med en lokal ring hjälte, går baren tyst. Malone vänder sig för att sehans fru, med ett ansikte dyster som död, förföljelse till baren.Slapping en fyra-bit bit ner på baren, drar hon sig upp till hennehela fem fot fem tum och säger till Mulcahey, "Ge mig vad själv harhar Havin alla dessa år. "Mulcahey tittar på Malone, som rycker på axlarna, och sedan tillbaka på Margaret MaryMalone. Han fastställer ett glas och häller henne en trippel skott av råg. Baren ärhelt tyst som de tittar på kvinnan plocka upp glaset och slå tillbakadryck. Hon slår glaset nedåt på stången, flämtar, ryser något ochsvimmar; falla rakt bakåt, stel som en styrelse, räddade från plötslig kontaktmed barroom golvet av riklig mage Seamus Fogerty.Någon gång senare, kommer hon att på bordet, en jacka under henneshuvud. Hennes blodsprängda ögon föll på hennes make, som säger: "Och alla dessaår du har thinkin "Jag har njutit meself."
		-- W. C. Fields, "My Little Chickadee"

%
Endast Irish coffee ger i ett enda glas alla fyra grundläggande matgrupper -alkohol, koffein, socker och fett.
		-- Alex Levine

%
Vänligen rök inte HÄR!Straff: En tidig, långsam död i cancer,emfysem, eller annan rökning-orsakad sjukdom.
		-- Alex Levine

%
Polisen: God kväll, är du värd?Värd: NejPolisen: Vi har fått klagomål om detta parti.Värd: Om drogerna?Polisen: Nej.Värd: Om vapnen, då? Är någon klagar vapnen?Polisen: Nej, buller.Värd: Åh, buller. Jo det är logiskt, eftersom det inte finns några vapeneller droger här. (En enorm explosion hörs ibakgrund.) Eller fyrverkerier. Vem klagar på buller?	Grannarna?Polisen: Nej, grannarna flydde inre timmar sedan. De flesta av de senasteklagomål har kommit från Pittsburgh. Tror du att du kundebe värd att lugna ner saker?Värd: No Problem. (Vid denna punkt, en Volkswagen bugg med primitivreligiösa symboler dras på dörrarna framgår av levanderum och ryter ner i korridoren, förbi polisen och pågräsmatta, där den slår i ett träd. Åtta gäster tumble utpå gräset, stönande.) Se? Saker och ting börjar att lindaner.
		-- Alex Levine

%
Syltdjurliv! En fest idag!
		-- Alex Levine

%
Recept för en Pan Galactic gurgla Blaster:(1) Ta saften från en flaska Ol 'Janx Spirit(2) Häll i det ett mått av vatten från havet avSantraginus V (Oh, de Santraginean fisk!)(3) Låt 3 kuber av Arcturan Mega-gin för att smälta in iBlandningen (korrekt iskallt eller bensin försvinner.)(4) Låt fyra liter Fallian kärr gas att bubbla genom den.(5) över baksidan av en silver sked, flyter ett mått påQualactin Hypermint extrakt.(6) Släpp i tanden av en Algolian Suntiger. Titta på den lösa.(7) Strö Zamphuor.(8) Lägg till en oliv.(9) Drinken ... men ... mycket noga ...
		-- Alex Levine

%
Riffle West Virginia är så liten att den scout fick fungera som denstad full.
		-- Alex Levine

%
Romantik, som alkohol, bör avnjutas, men bör inte tillåtas attbli nödvändig.
		-- Edgar Friedenberg

%
Sade den attraktiva, cigarr-rökare hemmafru till sin flickvän: "Jag fickbörjade en natt när George kom hem och fann en brinnande i askkoppen. "
		-- Edgar Friedenberg

%
Sam: Vad vet du det, Norm?Norm: Hur man sitta. Hur att dricka. Vill du frågesport mig?Sam: Hej, hur är livet behandlar dig där, Norm?Norm: Slår mig. ... Sen sparkar mig och lämnar mig att dö.Woody: Hur skulle en öl känner, mr Peterson?Norm: Ganska nervös om jag var i rummet.
		-- Cheers, Loverboyd

%
Sam: Vad är bra ord, Norm?Norm: Plop, plopp, fräsa, fräsa.Sam: Åh nej, inte den hungriga kviga ...Norm: Ja, ja, ja ...Sam: En halsbränna cocktail kommer upp.Sam: Whaddya säger Norm?Norm: Ja, jag har aldrig träffat en öl jag inte dricker. Och ner det går.Woody: Vad är din glädje, mr Peterson?Norm: Boxershorts och lösa skor. Men jag ska nöja sig med en öl.
		-- Cheers, The Bar Stoolie

%
Sam: Vad säger du, Norm?Norm: Alla billig, pråliga sak som får mig en öl.Sam: Vad säger du till en öl, Normie?Norm: Tjena, sjöman. Ny i stan?Norm: [kommer in från regnet] kväll, alla.All: normen! (Normand.)Sam: Fortfarande hälla Norm?Norm: Det är roligt, jag var på väg att be dig samma sak.
		-- Cheers, Diane's Nightmare

%
Sam: Vad är det som händer, Normie?Norm: Min födelsedag, Sammy. Ge mig en öl, hålla ett ljus i      det, och jag kommer att blåsa ut min lever.Woody: Hej, Mr P. Hur går sökandet efter Mr Calvin?Norm: Inte liksom sökandet efter Mr Donut.       Fann honom varje par av block.
		-- Cheers, Head Over Hill

%
Sam: Vad är nytt, Norm?Norm: De flesta av min fru.Coach: Öl, Norm?Norm: Naah, jag skulle förmodligen bara dricka det.Coach: Vad gör, Norm?Norm: Tja, vetenskap söker ett botemedel mot törst. jag råkar       vara marsvin.
		-- Cheers, Let Me Count the Ways

%
Visa respekt för ålder. Dricker gott Scotch för en förändring.
		-- Cheers, Let Me Count the Ways

%
Sömn - den mest vacker upplevelse i livet - utom dryck.
		-- W. C. Fields

%
Rökning är nu godkänd !!!Den som vill röka måste dock lämna, i tre exemplar, denUSA: s regering miljökonsekvensbeskrivning Narrative Statement (EINS)som i detalj beskriver den typ av förbränning som föreslås, påverkan påmiljö, och förväntade opposition. Uttalanden måste varainlämnad 30 dagar i förväg.
		-- W. C. Fields

%
Rökning är en av de främsta orsakerna till statistik.
		-- Fletcher Knebel

%
Rökning är, så vitt jag är orolig, hela poängen med att vara en vuxen.
		-- Fran Lebowitz

%
Rökning förbjuden. Absolut inga ifs, ands, eller rumpor.
		-- Fran Lebowitz

%
Så, är glaset halvtomt, halvfullt, eller bara dubbelt såstor som den behöver vara?
		-- Fran Lebowitz

%
Vissa människor har ingen respekt för ålder om det inte är på flaska.
		-- Fran Lebowitz

%
Ibland känner jag bara att hela världen är en cigarett och jag ärendast askkopp.
		-- Fran Lebowitz

%
Split 1/4 flaska .187 literHalv halv flaskaFlaska 750 milliliterMagnum 2 flaskor 1,5 literJeroboam 4 flaskorRehoboam 6 flaskor Ej tillgänglig i USAMethuselahs 8 flaskorSalmanazar 12 flaskorBalthazar 16 flaskorNebuchadnezzar 20 flaskor 15 literSovereign 34 flaskor 26 literThe Sovereign är en ny flaska, gjord för lanseringen avstörsta kryssningsfartyg i världen. Flaskan kostade 8000 dollaratt producera och de bara gjort åtta av dem.De flesta av de roliga namn kommer från bibliska personer.
		-- Fran Lebowitz

%
Symptom: Dricka inte ger smak och tillfredsställelse, är ölovanligt blek och klar.Problem: Glas tom.Nödvändiga åtgärder: Hitta någon som kommer att köpa dig en annan öl.Symptom: Dricka inte ger smak och tillfredsställelse,och framsidan av din skjorta är blöt.Fel: Mouth inte öppna när man dricker eller glas tillämpasfel del av ansiktet.Nödvändiga åtgärder: Köp en öl och praktik framför spegeln.Drick så många som behövs för att perfekt dricka teknik.
		-- Bar Troubleshooting

%
Symptom: Allt har gått mörkt.Fel: Bar stängs.Nödvändiga åtgärder: panik.Symptom: Du vaknar att hitta din säng hård, kall och våt.Du kan inte se badrum ljus.Fel: Du har tillbringat natten i rännstenen.Nödvändiga åtgärder: Kontrollera din klocka för att se om barer är öppna ännu. Om inte,Unna dig en lie-in.
		-- Bar Troubleshooting

%
Symptom: Fötterna kall och våt, glas tom.Fel: Glas hålls vid felaktig vinkel.Åtgärd krävs: Vrid glas på annat sätt så att öppna ändpunktermot taket.Symptom: fötter varma och fuktiga.Fel: Felaktig blåskontroll.Nödvändig åtgärd: Gå stå bredvid närmaste hund. Efter ett tag klagatill ägaren om sin brist på intern utbildning ochkräver en öl som kompensation.
		-- Bar Troubleshooting

%
Symptom: Golv suddig.Fel: Du bläddrar botten av tomma glas.Nödvändiga åtgärder: Hitta någon som kommer att köpa dig en annan öl.Symptom: Golv rörelse.Fel: Du genomförs.Nödvändig åtgärd: Ta reda på om du kommer till en annan bar. Om inte,klaga högljutt att du blir kidnappad.
		-- Bar Troubleshooting

%
Symptom: Golv gungande.Fel: Överdriven luftturbulens, kanske på grund av air-hockeyspel pågår.Åtgärd krävs: Sätt kvastskaftet ned baksidan av jackan.Symptom: Allt har gått svagt, konstig smak av jordnötteroch pretzels eller cigarettfimpar i munnen.Fel: Du har fallit framåt.Åtgärd krävs: Se ovan.Symptom: Motsatt vägg täckt med akustisk kakel och flerafluorescerande ljus remsor.Fel: Du har fallit bakåt.Nödvändiga åtgärder: Om glaset är fullt och ingen står pådricka arm, stanna kvar. Om inte, får någon att hjälpadu går upp, piska dig till bar.
		-- Bar Troubleshooting

%
Ta mig full, jag är hemma igen!
		-- Bar Troubleshooting

%
Det bästa publik är intelligent, välutbildad och lite berusad.
		-- Maurice Baring

%
Det bästa sättet att bevara en rätt är att utöva den, och rätten tillrök är en rätt värd att dö för.
		-- Maurice Baring

%
Kelterna uppfann två saker, whisky och självförstörelse.
		-- Maurice Baring

%
Kyrkan är nära men vägen är isig; baren är långt borta, men jag kommergå försiktigt.
		-- Russian Proverb

%
Levnadskostnaderna har just gått upp en annan dollar per liter.
		-- W. C. Fields

%
Fadern, som passerar genom sin sons college stad sent en kväll på enaffärsresa, trodde att han skulle betala sin pojke en suprise besök. Framme vidlad s broderskap hus, rapped pappa högt på dörren. Efter flera minuterknackar, drev en sömnig röst ned från en andra våningen fönster,"Whaddaya vill?""Gör Ramsey Duncan bor här?" frågade fadern."Ja", svarade rösten. "Dump honom på verandan."
		-- W. C. Fields

%
Ett tecken på en bra fest är att du vaknar upp nästa morgon villändra ditt namn och börja ett nytt liv i annan stad.
		-- Vance Bourjaily, "Esquire"

%
Sökandet efter den perfekta martini är ett bedrägeri. Den perfekta martini ärett bälte av gin från flaskan; något annat är de dekadenta grannlåtcivilisation.
		-- T.K.

%
Telefonen är ett bra sätt att prata med folk utan att behöva erbjudadem en drink.
		-- Fran Lebowitz, "Interview"

%
Domen av en jury är a priori yttrande som jurymedlem som rökerde värsta cigarrer.
		-- H. L. Mencken

%
Den yppiga blond chatta med hennes vackra eskort i en poshrestaurang när deras servitör, snubblande som han tog med sig sina drycker,dumpade en martini on the rocks ner på baksidan av den blonda klänning. Honsprang till hennes fötter med en vild rebell skrika, streckad vilt runt bordet,sedan galoppe wriggling från rummet följt av hennes distraught pojkvännen.En man som placeras på den andra sidan av rummet med ett datum av hans egna beckonedatt servitören och sade: "Vi kommer att ha två av vad hon drack."
		-- H. L. Mencken

%
Vattnet var inte passar att dricka. För att göra det tilltalande, vi var tvungna att lägga till whisky.Genom omsorgsfull ansträngning, lärde jag mig att gilla det.
		-- Winston Churchill

%
"Hela världen är cirka tre drinkar bakom."
		-- Humphrey Bogart

%
Den vise och intelligent kommer sent att inse att alkohol, ochinte hunden är människans bästa vän. Rover tar stryk - och han borde.
		-- W. C. Fields

%
Det finns fler gamla drinkare än gamla läkare.
		-- W. C. Fields

%
Det finns bara två typer av tequila. Bra och bättre.
		-- W. C. Fields

%
Det finns två problem med en stor baksmälla. Du kännersom du kommer att dö och du är rädd att du inte kommer.
		-- W. C. Fields

%
Det vara nyktra män a'plenty och drinkare knappt tjugo; det finns mänpå över nittio som har ännu aldrig kysst en flicka. Men ge mig vandringrover, från Orkney ner till Dover, kommer vi strövar omkring hela världen, ochtillsammans kommer vi att möta världen.
		-- Andy Stewart, "After the Hush"

%
Det är inget fel med avhållsamhet, med måtta.
		-- Andy Stewart, "After the Hush"

%
Det kommer alltid att finnas ölburkar rullar på golvet i bilen närchefen ber om skjuts hem från kontoret.
		-- Andy Stewart, "After the Hush"

%
Dessa dagar livets nödvändigheter kostar ungefär tre gånger mer än vad devan vid, och halva tiden är de inte ens passar att dricka.
		-- Andy Stewart, "After the Hush"

%
De tog några av Van Goghs, de flesta av juvelerna, och alla Chivas!
		-- Andy Stewart, "After the Hush"

%
Att vara berusad är att känna sofistikerad men inte kunna säga det.
		-- Andy Stewart, "After the Hush"

%
Till en stor kalkon lägga en gallon vermouth och en damejeanne av Angosturabitter. Skaka.
		-- F. Scott Fitzgerald, recipe for turkey cocktail.

%
Alltför slet. Måste gå.
		-- F. Scott Fitzgerald, recipe for turkey cocktail.

%
Tandkräm skadar aldrig smaken av god whisky.
		-- F. Scott Fitzgerald, recipe for turkey cocktail.

%
Två vänner var ute dricka när plötsligt en krängde bakåt av sigbarstol och låg orörlig på golvet."En sak om Jim," den andra sa till bartendern, "han säkervet när du ska sluta. "
		-- F. Scott Fitzgerald, recipe for turkey cocktail.

%
Vermouth gör mig alltid lysande om det gör mig idiotiskt.
		-- E. F. Benson

%
Vi röker inte och vi inte tugga, och vi inte gå med tjejer som gör det.
		-- Walter Summers

%
Vilken skurk stal korken ur min lunch?
		-- J. D. Farley

%
När allt annat misslyckas, häll en pint Guinness i bensintanken, avanceratänd 20 grader, gråta "God Save the Queen", och dra i startvredet.
		-- MG "Series MGA" Workshop Manual

%
När jag dricker, "en man ropade * allas * drycker till de församlade bar mecenater.Ett högt allmänt jubel gick upp. Efter Downing sin whisky, hoppade han på enbarstol och ropade "När jag tar en drink, * alla * tar en annandricka! "Tillkännagivandet producerade en annan glädje och en annan runda av drycker.Så snart han hade downed sin andra drink, hoppade stipendiaten tillbakapå pallen. "Och när jag betalar" han vrålade, slapping fem dollar påbaren "* alla * lönar sig!"
		-- MG "Series MGA" Workshop Manual

%
När jag värms mitt hem med olja, använde jag i genomsnitt 800 liter per år. jaghar funnit att jag kan hålla bekvämt varma för en hel vinter meddrygt hälften mängd öl.
		-- Dave Barry, "Postpetroleum Guzzler"

%
När jag säljer sprit, det kallas bootlegging; när mina patrons tjänardet på silverbrickor på Lake Shore Drive, det kallas gästfrihet.
		-- Al Capone

%
När koppen är full, bära den nivå.
		-- Al Capone

%
När det blir tufft, den tuffa gå ta en öl.
		-- Al Capone

%
Medan ridning i ett tåg mellan London och Birmingham, en kvinnafrågade Oscar Wilde: "Du har inget emot om jag röker, eller hur?"Wilde gav henne en sidoblick och svarade: "Jag har inget emot omdu bränner, fru. "
		-- Al Capone

%
Vem behöver vänner, när du kan sitta ensam i rummet och dricker?
		-- Al Capone

%
Varför i hela friden gör folk köper gamla flaskor vin när de kan få enfärskt för en fjärdedel av priset?
		-- Al Capone

%
Kvinna på gatan: Sir, du är full; mycket, mycket berusade.Winston Churchill: Madame, är du ful; mycket, mycket ful.Jag ska vara nykter på morgonen.
		-- Al Capone

%
Underbar dag. Din baksmälla gör bara det verkar fruktansvärt.
		-- Al Capone

%
Woody: Vad är historien, mr Peterson?Norm: De Bobbsey tvillingar gå till bryggeriet.        Låt oss bara klippa till det lyckliga slutet.Woody: Hej, mr Peterson, finns det en kall väntar på dig.Norm: Jag vet, och om hon ringer, jag är inte här.Sam: Öl, Norm?Norm: Har jag fått det förutsägbara? Bra.
		-- Cheers, Don't Paint Your Chickens

%
Woody: Hej, mr Peterson, Jack Frost löste på näsan?Norm: Japp, nu ska vi få Joe öl löste på min lever, va?Sam: Vad är du upp till Norm?Norm: Min idealvikt om jag var elva fot lång.Woody: Nice kall öl kommer upp, mr Peterson.Norm: Du menar, `trevlig kall öl går * ner * Mr Peterson.
		-- Cheers, Loverboyd

%
Woody: Hej, mr Peterson, vad säger du till en kall?Norm: Vi ses senare, Vera, jag ska vara på Cheers.Sam: Tja, titta på dig. Du ser ut som katten som svalde kanariefågeln.Norm: Och jag behöver en öl att skölja ner honom.Woody: Vill du ha en öl, mr Peterson?Norm: Nej, jag vill ha en död katt i ett glas.
		-- Cheers, Little Carla, Happy at Last, Part 2

%
Woody: Hej, vad är mr Peterson upp?Norm: Garantin på min lever.Sam: Vad kan jag göra för dig, Norm?Norm: Öppna upp dessa öl kranar och, oh, ta ledigt, Sam.Woody: Vad som händer, mr Peterson?Norm: Ett annat skikt för vintern, trä.
		-- Cheers, It's a Wonderful Wife

%
Woody: Hur mår du idag, Mr. Peterson?Norm: Dålig.Woody: Åh, jag är ledsen att höra det.Norm: Nej, jag menade 'pour'.Woody: Hej, vad är Mr Peterson historien?Norm: Boy meets öl. Pojke dricker öl. Pojke får en annan öl.Paul: Hej Norm, hur världen behandlat dig?Norm: Som ett barn behandlar en blöja.
		-- Cheers, Tan 'n Wash

%
Woody: Vad som händer, mr Peterson?Norm: Låt oss tala om vad som händer * i * Mr Peterson. En öl, Woody.Sam: Hur liv behandlar dig?Norm: Det är inte, Sammy, men det betyder inte att du inte kan.Woody: Kan jag häller dig ett förslag, mr Peterson?Norm: En lite tidigt, är det inte Woody?Woody: För en öl?Norm: Nej, för dumma frågor.
		-- Cheers, Let Sleeping Drakes Lie

%
Woody: Vad händer, mr Peterson?Norm: Frågan är, Woody, varför är det som händer med mig?Woody: Vad händer ner, mr Peterson?Norm: Mina kinder på denna barstol.Woody: Hej, Mr Peterson kan jag hälla en öl?Norm: Ja, okej, Woody, men tänk på att stoppa mig på en. ...       Eh, göra det 1-30.
		-- Cheers, Strange Bedfellows, Part 2

%
Arbete är förbannelsen av dricka klasser.
		-- Mike Romanoff

%
Du kan inte falla från golvet.
		-- Mike Romanoff

%
Du är inte en alkoholist om du går till mötena.
		-- Mike Romanoff

%
Du är inte druckit om du kan ligga på golvet utan att hålla på.
		-- Dean Martin

%
