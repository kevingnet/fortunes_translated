En viss gammal katt hade gjort sitt hem i gränden bakom Gabe bar för vissatid, lever på rester och enstaka stenciler från bartendern. Enkväll, uppmuntrat av hunger, kattdjur försökte följa Gabe genombakdörren. Tyvärr hade bara hans kropp tagit sig igenom närdörren stängdes, bryta kattens svans vid sin bas. Detta visade sig vara alltförmycket för den gamla varelse, som såg sorgset på Gabe och löpte på plats.Gabe sätta stommen tillbaka ut i gränden och gick tillbaka till verksamheten.Den obligatoriska stängningstid kom och Gabe var i färd med att låsa uppefter de sista kunderna hade gått. Närmar bakdörren han blev överraskadatt se en uppenbarelse av det gamla katt mournfully hålla sitt avhuggna svans ut,tyst pläderar för Gabe att sätta svans tillbaka på sin kropp så att den kundegå vidare till kitty after komplett.Gabe skakade sorgset på huvudet och sade till spöke, "jag kan inte. Du vetlagen - ingen detaljhandel sprit efter 02:00 ".
		-- Will Rogers

%
En landsman mellan två advokater är som en fisk mellan två katter.
		-- Ben Franklin

%
En läkare var strandsatta med en advokat i en läckande livflotte i haj-smittadevattnen. Läkaren försökte simma i land men åts av hajar. Deadvokat, dock simmade säkert förbi blodtörstiga hajar. "Professionellartighet ", förklarade han.
		-- Ben Franklin

%
A Dublin advokat dog i fattigdom och många advokater i staden prenumererar påen fond för hans begravning. Den Lord Chief Justice Orbury ombads att doneraen shilling. "Bara en shilling?" utbrast mannen. "Endast en shilling att begravaen advokat? Här är en försöks; gå och begrava tjugo av dem. "
		-- Ben Franklin

%
En vän till mig kommer inte att få en skilsmässa, eftersom han hatar advokater mer än hanhatar hans hustru.
		-- Ben Franklin

%
En grundskola lärare frågade eleverna vad deras föräldrar gjordeför ett levande. "Tim, du först", sade hon. "Vad gör din mamma görahela dagen?"Tim stod upp och stolt sa: "Hon är en läkare.""Det är underbart. Vad säger du, Amie?"Amie blygt stod upp, scuffed hennes fötter och sade: "Min far är enbrevbärare.""Tack, Amie," sa läraren. "Och din far, Billy?"Billy stod stolt upp och meddelade, "Min pappa spelar piano i enhorhus."Läraren var bestört och snabbt bytte till geografi.Senare samma dag gick hon till Billys hus och ringde. Billys pappasvarade dörren. Läraren förklarade vad hans son hade sagt och krävten förklaring.Billys far svarade: "Ja, jag är verkligen en advokat. Men hur gördu förklara något sådant till ett sju år gammalt barn? "
		-- Ben Franklin

%
En hemmafru, en revisor och en advokat ombads att lägga två och två.Husmodern svarade: "Four".Revisorn sade, "Det är antingen 3 eller 4. Låt mig köra dessa siffrorgenom min kalkylbladet en gång. "Advokaten drog draperier, nedtonade ljus och bad i endämpad röst, "Hur mycket vill du att det ska vara?"
		-- Ben Franklin

%
En jury består av tolv personer valt att avgöra vem som har bättre advokat.
		-- Robert Frost

%
En advokat som heter Strange var shopping för en gravsten. Efter han hadegjort sitt val, frågade stenhuggare honom vad inskrift hanvill på det. "Här ligger en ärlig man och en advokat," svaradeadvokat."Tyvärr, men jag kan inte göra det", svarade stenhuggare. "I dennatillstånd, är det mot lagen att begrava två personer i samma grav. Dock,Jag skulle kunna sätta `` här ligger en ärlig advokat ', om det skulle vara okej. ""Men det kommer inte att låta folk veta vem det är" protesterade advokaten."Visst kommer", svarade den stenhuggare. "Människor kommer att läsa detoch utropa: "Det är märkligt!"
		-- Robert Frost

%
En Los Angeles domare ansåg att "en medborgare kan snarka med immunitetsitt eget hem, även om han kan vara i besittning av ovanlig ochexceptionella förmåga att visst område. "
		-- Robert Frost

%
En Los Angeles domare ansåg att "en medborgare kan snarka med immunitetsitt eget hem, även om han kan vara i besittning av ovanliga och exceptionellaförmåga att visst område. "
		-- Robert Frost

%
En man gick in i en bar med sin alligator och frågade bartendern,"Vill du tjäna advokater här?"."Visst gör", svarade bartendern."Bra", sa mannen. "Ge mig en öl, och jag kommer att ha en advokat förmin "gator".
		-- Robert Frost

%
A New York domare slagit fast att om två kvinnor bakom dig påfilmer insisterar på att diskutera den sannolika resultatet av filmen, har durätt att vända och blåsa en Bronx jubel på dem.
		-- Robert Frost

%
A New York förordningen förbjuder inspelningen av kaniner frånbaksida en Third Avenue gata bil - om bilen är i rörelse.
		-- Robert Frost

%
En Riverside, Kalifornien, hälsa förordningen sägs att två personer kaninte kyssa varandra utan att först torka sina läppar med carbolized rosenvatten.
		-- Robert Frost

%
En liten stad som inte kan stödja en advokat kan alltid att stödja två.
		-- Robert Frost

%
Enligt Arkansas lag, avsnitt 4761, påvens Digest: "Ingen personskall tillåtas under någon förevändning som helst, för att komma närmare änfemtio fot av någon dörr eller ett fönster av någon röstningen rum, från öppningenav röstningarna fram till slutförandet av räkningen och certifiering avavkastningen. "
		-- Robert Frost

%
Enligt Kentucky nationell lag, måste varje person ta ett bad åtminstoneen gång om året.
		-- Robert Frost

%
Efter 35 år, har jag avslutat en omfattande studie av den europeiskakomparativ rätt. I Tyskland, enligt lagen, är allt förbjudet,utom det som är tillåtet. I Frankrike, enligt lag, alltär tillåtet, utom det som är förbjudet. I Sovjetunionen,enligt lagen, är allt förbjudet, inklusive det som ärtillåten. Och i Italien, enligt lagen, allt är tillåtet,särskilt det som är förbjudet.Tal till Association of American Law skolor, 1985
		-- Newton Minow,

%
Efter hans Ignoble Disgrace, Satan höll på att utvisas frånHimmel. När han passerade genom grindarna, stannade han ett ögonblick i tanken,och vände sig till Gud och sa: "En ny skapelse kallad Man, jag hör, är snartsom ska skapas. ""Detta är sant", svarade han."Han kommer att behöva lagar", sade Demon slugt."Vad! Du, den bestämda Enemy för all framtid! Du ber om deträtt att göra sina lagar? "	"Å nej!" Satan svarade: "Jag ber bara att han tillåtas attgöra sin egen. "Det var så beviljades.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
En ändring av en rörelse kan ändras, men en ändring till en ändringtill en rörelse som inte kan ändras. Men ett substitut för en ändring avoch ändring av en rörelse kan antas och ersättaren kan ändras.språk.
		-- The Montana legislature's contribution to the English

%
En advokat försvarade sin klient mot en avgift på mord."Your Honor är min klient anklagas för fyllning sin älskares stympade kropp ien resväska och på väg till den mexikanska gränsen. Strax norr om Tijuana en polisfläckig handen sticker ut ur resväskan. Nu, jag vill betonaatt min klient är * ___ inte * en mördare. En slarvig packare, kanske ... "
		-- The Montana legislature's contribution to the English

%
En engelsk domare, växande trötta på advokatlångrandig summering,lutade sig över bänken och sade: "Jag har hört era argument, SirGeoffrey och jag är klokare! "Sir Geoffrey svarade:" Det kan vara,Milord, men åtminstone du är bättre informerade! "
		-- The Montana legislature's contribution to the English

%
Och så var det advokat som ingrep kogödsel och tankehan smälte ...
		-- The Montana legislature's contribution to the English

%
En annan dag, en annan dollar.på Hinckleys frikännande för fotografering president RonaldReagan.
		-- Vincent J. Fuller, defense lawyer for John Hinckley,

%
Antitrustlagar bör behandlas med exakt den attityden.
		-- Vincent J. Fuller, defense lawyer for John Hinckley,

%
Atlanta gör det olagligt att knyta en giraff till en telefonstolpeeller gatlykta.
		-- Vincent J. Fuller, defense lawyer for John Hinckley,

%
Justitiekansler Edwin Meese III förklarade varför Högsta domstolens Mirandabeslut (innehav att patienter har rätt att tiga och har enadvokat närvarande vid förhör) är onödig: "Du har inte mångamisstänkta som är oskyldig för ett brott. Det är motsägelsefullt. Om en personär oskyldig till brott, då är han inte en misstänkt. "
		-- U.S. News and World Report, 10/14/85

%
Var uppriktig och tydlig med din advokat ... är det hans sak att förvirrafrågan efteråt.
		-- U.S. News and World Report, 10/14/85

%
Se garantin - det fetstil giver och finstilta tager bort.
		-- U.S. News and World Report, 10/14/85

%
Att vara en gruvarbetare, så fort du är för gammal och trött och sjuk och dumt attgör ditt jobb ordentligt, måste du gå, där det motsatta gäller meddomarna.
		-- Beyond the Fringe

%
Mellan grand theft och en rättslig avgift, bara det står en juristexamen.
		-- Beyond the Fringe

%
... Men som register över domstolar och rättvisa är tillåtlig, det kan lätt varavisat att kraftfulla och illvilliga trollkarlar gång fanns och var ett gisselmänskligheten. Bevisen (inklusive bekännelse) vid vilken vissa kvinnordömdes för häxeri och avrättades var utan fel; det är fortfarandeoförvitlig. Domarnas beslut baserade på det var ljud i logik ochi lagen. Ingenting i befintliga domstol någonsin mer noggrant bevisat änanklagelserna om häxkonst och trolldom som så många led döden. Omdet fanns inga häxor, mänsklig vittnesbörd och mänskligt förnuft är likadana utblottadeav värde.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Carmel, New York, har en förordning som förbjuder män att bära rockar ochbyxor som inte matchar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Vissa passager i flera lagar har alltid trotsat tolkning ochmest oförklarlig måste vara en bedömningsfråga. En domare av revisionsSession of Scotland har sänt redaktörerna för boken hans kandidat somlyder: "I Nuts (oslipade), (andra än jordnötter) Order, uttrycketnötter skall ha hänvisning till sådana nötter, andra än jordnötter, som skullemen för denna ändrings Order inte som nötter (oslipade) (andra än markmuttrar) på grund av att de är nötter (oslipade). "
		-- Guiness Book of World Records, 1973

%
Chicago lag förbjuder äta på en plats som är på brand.
		-- Guiness Book of World Records, 1973

%
Diogenes gick för att leta efter en ärlig advokat. "Hur går det?", Någonfrågade honom efter några dagar."Not too bad", svarade Diogenes. "Jag har fortfarande min lykta."
		-- Guiness Book of World Records, 1973

%
[District Advokatbyrå] lära i District Attorney skolan att det finnstvå bergsäkert sätt att få en hel del positivt publicitet:(1) Gå ner och raid alla skåp i den lokala high school och    konfiskera 53 marijuanacigaretter och lägg dem i en hög och håll    en presskonferens där man tillkännager att de har ett värde på gatan    av $ 850.000.000. Dessa räder aldrig misslyckas, eftersom alla högstadier,    inklusive helt nya, aldrig använda dem, har åtminstone 53 marijuana    cigaretter i skåpen. Såvitt någon kan berätta, locker    Fabriken sätter dem där.(2) Raid en "vuxen bok butik" och hålla en presskonferens där man    meddelar du laddar ägare med 850 punkter för att vara en    bit av human sleaze. Detta också misslyckas aldrig, eftersom du alltid    få en fällande dom. En jurymedlem vid en pornografi rättegången handlar inte om att    tillstånd för den post som han finner inget obscent om en film    där aktörer delta i sexuella aktiviteter med levande ormar och en    brandsläckare. Han kommer att döma bokhandeln ägare, och    rösta för dödsstraffet bara för att se till att ingen blir fel    intryck.
		-- Dave Barry, "Pornography"

%
District of Columbia fotgängare som hoppar över passerande bilar att flyskada, och sedan slå bilen när de kommer ner, är ansvarig för eventuellaskadorna på fordonet.
		-- Dave Barry, "Pornography"

%
Skilsmässa är ett spel som spelas av advokater.
		-- Cary Grant

%
Läkare och advokater måste gå till skolan år efter år, ofta medlite sömn och med stor uppoffring för sina första fruar.
		-- Roy G. Blount, Jr.

%
Slagsmål mellan katter och hundar är förbjudna enligt lag i Barber, NorthCarolina.
		-- Roy G. Blount, Jr.

%
Först var Dial-A-bön, sedan Dial-A-recept, och även Dial-A-fotbollsspelare.Men sydöstra viktorianska staden Sale har producerat en till toppen dem alla.Dial-A-Wombat.Det hela började tidigt igår när Sale polisen fick ett telefonsamtalring: "Du kommer inte tro det, och jag är inte full, men det finns en wombat itelefonkiosk utanför stadshuset ", den som ringer säger.Inte övertygad om om den som ringer anspråk på nykterhet, medlemmar iden Constabulary körde till platsen, räknar med att plocka upp en berusad.Men där var det en irriterad wombat, instängd i en telefonkiosk.Den wombat, fast besluten att inte vara hade det bättre av igen, kastade sinbulk in i striden. Det var slutligen lassoed och släpptes i en närliggande scrub.Sedan fick officerarna annat meddelande ... en annan wombat ien annan telefonkiosk.Det var det: * En annan * arg wombat instängd i en telefonkiosk.Konstaplarna tog miffed pungdjur i tillfälligt förvar ochsläppt det, även i skurar.Men på väg tillbaka till stationen de råkade passera en annantelefonkiosk, och - du gissade det - en annan fängslade wombat.Efter några allvarliga detektivarbete, grabbarna i blått hittat en misstänkt,och efter förhör, släppte honom som tas ut på kallelsen.Deras problem ... de kan inte hitta en lag mot att placera wombats itelefonkiosker.
		-- "Newcastle Morning Herald", NSW Australia, Aug 1980.

%
För vissa människor, efter femtio, tar tvister platsen för kön.
		-- Gore Vidal

%
För tre år hade den unge advokat tagit hans kortsemester på detta land inn. Sista gången han hade äntligen enaffär med gästgivare dotter. Ser fram emot en spännandenågra dagar, drog han sin resväska uppför trapporna av inn, sedan slutadekort. Där satt sin älskare med ett spädbarn på knät!"Helen, varför inte du skriver när du lärt du var gravid?"han grät. "Jag skulle ha rusat upp här, vi kunde ha gift,och barnet skulle ha mitt namn! ""Jo", sa hon, "när mina föräldrar fick reda på mitt tillstånd,Vi satt uppe hela natten pratar och pratar och slutligen bestämde att det skulle varabättre att ha en jävel i familjen än en advokat. "
		-- Gore Vidal

%
Fortune dokumenterar stora rättsliga beslut:Det är en bevisregel härledas från upplevelsen av mänskligheten ochstöds av förnuft och myndighet som positiva vittnesbörd har rätt tillmer vikt än negativa vittnesmål, men den senare termen menasnegativ vittnesbörd i dess rätta bemärkelse och inte bevis på ennegativt, eftersom vittnesbörd till stöd för en negativ kan vara så positivsom stöd för ett jakande.
		-- 254 Pac. Rep. 472.

%
Fortune dokumenterar stora rättsliga beslut:Vi kan föreställa oss ingen anledning, med vanlig omsorg, kunde mänskliga tårna inte varautelämnats av tuggtobak, och om tårna finns i tuggtobak, detverkar för oss att någon har varit mycket oförsiktig.
		-- 78 So. 365.

%
Fortune dokumenterar stora rättsliga beslut:Vi tror att vi kan ta rättsliga meddelande om att begreppet "bitch"kan innebära en viss känsla av smekning när den tillämpas på en kvinna i hundart men att det är sällan, om någonsin, så används när det tillämpas på en kvinnligav den mänskliga rasen. Kommer som det gjorde, ganska nära i hälarna på tvårevolverskott riktade mot personen som det användes troligen, vi trordet bär varje rimlig konsekvens av illvilja mot den personen.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortune lag av veckan (den här veckan, från Kentucky):Ingen kvinna ska visas i en baddräkt på någon flygplats i dettaStat, såvida hon eskorteras av två tjänstemän eller om hon är beväpnadmed en klubb. Bestämmelserna i denna stadga skall inte tillämpas på kvinnorväger mindre än 90 pounds eller mer än 200 pounds, inte heller skall dettillämpas på kvinnliga hästar.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortune utnämning för All-Time mästare och beskyddare av ungdomligMoral går till representant Clare E. Hoffman of Michigan. under enpassionerad House debatten om ett lagförslag för att "expandera ostron ochclam forskning ", en skarp öron informant transkriberas följandeutbyte mellan vår hjälte och tekniker. John D. Dingell, även Michigan.Dingell: Det finns platser i världen i dagsläget där vi ärbehöva artificiellt propagera ostron och musslor.HOFFMAN: Du menar ostron jag köper inte naturens ostron?Dingell: De kan eller inte kan vara naturlig. Det enkla faktumär att kvinnliga ostron genom sina levnadsvanor kasta utstora mängder utsäde och de manliga ostron kastade ut storamängder av gödsling ...HOFFMAN: Vänta en minut! Jag vill inte gå in på det. Det är mångatonåringar som läser Congressional Record.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 18:Q: Är du gift?A: Nej, jag är frånskild.Fråga: Och vad gjorde din man göra innan du frånskild honom?A: En hel del saker som jag inte visste om.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 19:Fråga: Doktorn, hur många obduktioner har du utfört på döda människor?A: Alla mina obduktioner har utförts på döda människor.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 25:F: Du säger att du hade tre män stans på dig, sparka dig, våldta dig,    och du inte skrika?S: Nej frun.F: Betyder att du samtyckt?A: Nej, frun. Det innebär att jag var medvetslös.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 29:DOMAREN: Nu när vi börjar, måste jag be er att bannlysa alla närvarandeInformation och fördomar från dina sinnen, om du har någon ...
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 32:Q: Vet du hur långt gravid du är just nu?A: Jag kommer att vara tre månader 8 november.Q: Tydligen sedan, dagen för befruktningen var 8 augusti?A: Ja.Fråga: Vad gjorde du och din man gör på den tiden?
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 37:Fråga: Har han plocka hunden upp i öronen?A: Nej.F: Vad gjorde han med hundens öron?A: Plocka upp dem i luften.F: Var var hunden vid den här tiden?A: I anslutning till öronen.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal citat # 3:F: När han gick, hade du gått och hon hade, om hon ville och var    stånd, för närvarande med undantag för alla begränsningar på henne att inte    gå, borta också, skulle han ha fört dig, vilket innebär att du och hon, med    honom till stationen?HERR. BROOKS: invändning. Frågan bör tas ut och sköt.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 41:Fråga: Nu, Mrs. Johnson, hur var din första äktenskap avslutas?A: Genom döden.Q: Och vars död den avslutade?
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal Citat # 52:F: Vad är ditt namn?A: Ernestine McDowell.F: Och vad är ditt civilstånd?En marknad.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Fortunes verkliga livet rättssal citat # 7:Fråga: Vad hände då?A: Han berättade, säger han, "Jag måste döda dig eftersom du kan identifiera mig."Fråga: Har han döda dig?A: Nej.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Frankfort, Kentucky, gör det olagligt att skjuta ut en polis tie.
		-- Smith v. Moran, 193 N.E. 2d 466.

%
"Gentlemen av juryn,", sade försvarsadvokat, börjar nuvärmas upp till sin summering ", den verkliga frågan här innan du är, skall dettavacker ung kvinna tvingas att tyna bort bort sina vackraste år i enmörk fängelsecell? Eller skall hon bli fria att återvända till sin mysiga lillalägenhet på 4134 Mountain Ave. - Där för att tillbringa sin ensamma, loveless timmari sin boudoir, liggande bredvid sin lilla prinsessa telefon, 962-7873? "
		-- Smith v. Moran, 193 N.E. 2d 466.

%
Komma sparkas ut ur American Bar Association är omtyckt få sparkasur boken-of-the-Month Club.av American Bar Association
		-- Melvin Belli on the occcasion of his getting kicked out

%
Gud bestämde sig för att ta djävulen till domstol och lösa sina meningsskiljaktigheteren gång för alla.När Satan hörde detta, flinade han och sa, "Och just där nitror du kommer att hitta en advokat? "
		-- Melvin Belli on the occcasion of his getting kicked out

%
Bra regeringen beror aldrig på lagar, men på de personliga egenskaperde som styr. Maskineri regeringen är alltid underordnadkommer av dem som administrerar det maskiner. Den viktigaste delen avregering, därför, är metoden för att välja ledare.
		-- Frank Herbert, "Children of Dune"

%
Han är ingen advokat som inte kan ta två sidor.
		-- Frank Herbert, "Children of Dune"

%
"Hej, jag heter Preston A. Mantis, vd för konsumenter Retail lag Outlet. Som nikan se genom min kostym och det faktum att jag har alla dessa böcker av samma höjdpå hyllorna bakom mig, jag är utbildad laglig advokat. Har du en bileller ett jobb? Har du någonsin gå runt? Om så är fallet, har du förmodligen ärendes aven utmärkt rättsfall. Även om det naturligtvis varje fall är olika, jagskulle definitivt säga att utifrån min erfarenhet och utbildning, det finns ingenanledningen till att du inte bör komma ut ur den här saken med åtminstone en stugakryssare."Kom ihåg, i Preston A. Mantis Konsumenter Retail lag Outlet, vårt mottoär: "Det är mycket svårt att motbevisa vissa typer av smärta."
		-- Dave Barry, "Pain and Suffering"

%
Hästar är förbjudet att äta brandposter i Marshalltown, Iowa.
		-- Dave Barry, "Pain and Suffering"

%
How do you förolämpa en advokat?Du kan lika gärna inte ens försöka. Överväg: av alla starktutbildad och utbildade yrken, är lagen den enda där det främstalärdom är att * vinna * är viktigare än * sanning *.När någon har sjunkit till den nivån, vad värre kan du säga om dem?
		-- Dave Barry, "Pain and Suffering"

%
HR 3128. Omnibus Budget Reconciliation, Fiscal 1986. Martin, R-Ill., Rörelseatt huset avta från sin oenighet till senaten ändringen görförändringar i propositionen att minska skatte 1986 underskott. Senaten ändringvar en ändring till kammaren ändring av senaten ändring av kammarenändring av senaten ändring av räkningen. Den ursprungliga Senate ändringvar konferensavtalet på räkningen. Enats om att.
		-- Albuquerque Journal

%
Humor i th domstolen:Fråga: Dricker du när du är i tjänst?A: Jag dricker inte när jag är i tjänst, om jag kommer på tull berusad.
		-- Albuquerque Journal

%
Humor i domstolen:Q. Och slutligen, Gary, måste alla dina svar vara muntligt. OK.? Vilken skola göra    du går till?A. Oral.Fråga: Hur gammal är du?A. Oral.
		-- Albuquerque Journal

%
Humor i domstolen:F. Och vem är denna person du talar om?A. Min ex-änka sa det.
		-- Albuquerque Journal

%
Humor i domstolen:F. Har du någonsin stanna hela natten med denna man i New York?A. Jag vägrar att svara på den frågan.F. Har du någonsin stanna hela natten med den här mannen i Chicago?A. Jag vägrar att svara på den frågan.F. Har du någonsin stanna hela natten med den här mannen i Miami?S. Nej
		-- Albuquerque Journal

%
Humor i domstolen:Q. Doktor, sa du att han blev skjuten i skogen?S. Nej, sa jag att han blev skjuten i ländryggen.
		-- Albuquerque Journal

%
Humor i domstolen:Q. Mrs Jones, är ditt utseende i morse i enlighet med en avsättning    märker som jag skickade till din advokat?S. Nej Detta är hur jag klär när jag går till jobbet.
		-- Albuquerque Journal

%
Humor i domstolen:Q. Mrs Smith, tror du att du är känslomässigt instabil?A. Jag borde vara.Fråga: Hur många gånger har du begick självmord?A. Fyra gånger.
		-- Albuquerque Journal

%
Humor i domstolen:Q. Officer, vad som ledde dig att tro att svaranden var påverkad?A. Eftersom han var argumentary och han kunde inte pronunciate hans ord.
		-- Albuquerque Journal

%
Humor i domstolen:F. Var du förtrogen med den avlidne?A. Ja, sir.F. Före eller efter hans död?
		-- Albuquerque Journal

%
Humor i domstolen:Fråga: Vad är din bror-i-lags namn?A. Borofkin.Fråga: Vad är hans förnamn?A. Jag kan inte minnas.Q. Han har varit din bror-in-law för år, och du kan inte komma ihåg sin första    namn?A. Nej, jag säga att jag är alltför upphetsad. (Resning från vittnesstolen och    pekar på Mr Borofkin.) Nathan, för Guds skull, berätta din första    namn!
		-- Albuquerque Journal

%
Humor i domstolen:Q: (Visar man bilden.) Det är du?A: Ja, sir.Q: Och du var närvarande när bilden togs, eller hur?
		-- Albuquerque Journal

%
Humor i domstolen:Q: ... och vad gjorde han då?A: Han kom hem, och nästa morgon var han död.Q: Så när han vaknade upp nästa morgon var han död?
		-- Albuquerque Journal

%
Humor i domstolen:Q: ... några förslag på vad hindrade detta från att vara en mordrättegång   i stället för ett försök till mordrättegång?A: Offret levde.
		-- Albuquerque Journal

%
Humor i domstolen:Q: Är du kvalificerad att ge ett urinprov?A: Ja, jag har varit sedan tidig barndom.
		-- Albuquerque Journal

%
Humor i domstolen:Q: Är du sexuellt aktiv?A: Nej, jag ligger bara där.
		-- Albuquerque Journal

%
Humor i domstolen:Fråga: Kan du se honom från där du stod?A: Jag kunde se hans huvud.Q: Och där var hans huvud?A: Precis ovanför axlarna.
		-- Albuquerque Journal

%
Humor i domstolen:Fråga: Har du berätta din advokat att din man hade erbjudit dig kränkningar?A: Han ville inte ge mig ingenting; han bara sa att jag kunde ha möbler.
		-- Albuquerque Journal

%
Humor i domstolen:Q: Nu har du undersökt andra mord, har du inte, där det fanns   ett offer?
		-- Albuquerque Journal

%
Humor i domstolen:Fråga: Så, efter bedövning, när du kom ut ur det, vad gjorde du observerar   med avseende på hårbotten?A: Jag såg inte min hårbotten hela tiden jag var på sjukhuset.Fråga: Det var täckt?A: Ja, bandagerade.Fråga: Sedan, senare .. vad såg du?A: Jag hade en hudtransplantation. Hela min skinkor och ben togs bort och sätta på toppen   mitt huvud.
		-- Albuquerque Journal

%
Humor i domstolen:F: Sanningen är att du inte var en opartisk, objektiv   vittne, är det inte. Du var alltför skjuten i bråken?A: Nej, sir. Jag blev skjuten halvvägs mellan bråken och örlogsfartyg.
		-- Albuquerque Journal

%
Humor i domstolen:Q: Vad kan du berätta om sanningshalten och sanningshalten i denna svarande?A: Åh, hon kommer att berätta sanningen. Hon sade att hon skulle döda den sonofabitch - och   hon gjorde!
		-- Albuquerque Journal

%
Humor i domstolen:Fråga: Vad är innebörden av spermier är närvarande?A: Det indikerar samlag.Q: Man spermier?A. Det är den enda sorten jag vet.
		-- Albuquerque Journal

%
Humor i domstolen:Fråga: Vilket är ditt förhållande med käranden?A: Hon är min dotter.Q: Var hon din dotter på 13 Februari 1979?
		-- Albuquerque Journal

%
Jag behöver en annan advokat som jag behöver ett annat hål i mitt huvud.
		-- Fratianno

%
Jag minns när laglig används för att betyda laglig, nu det innebär någratyp av lucka.
		-- Leo Kessler

%
Jag antar att en del av variationen mellan Boston förare och resten avland beror på den progressiva Massachusetts förarutbildning Manual somJag råkar ha i min topp skrivbordslåda. Några av de tips för bättre körningär värt att överväga, nämligen:[110,13]:       "När du reser på en enkelriktad gata, stanna till höger, så att inte        störa mötande trafik. "[22.17b]:       "Att lära sig att byta fil tar tid och tålamod. Det bästa        rekommendation som kan göras är att gå till en Celtics [basket]        spel; studera snabb paus och sedan gå ut och praktisera det        på motorvägen. "[41,16]:       "Bump aldrig en barnvagn av ett övergångsställe om barnet är verkligen        ber om det."
		-- Leo Kessler

%
Jag antar att en del av variationen mellan Boston förare och resten avland beror på den progressiva Massachusetts förarutbildning Manual somJag råkar ha i min topp skrivbordslåda. Några av de tips för bättre körningär värt att överväga, nämligen:[131.16d]:       "Körriktningsvisare i allmänhet inte används förutom under fordonet        inspektion; emellertid är en vänster-sväng signal lämplig när man gör        en U-sväng på en delad highway. "[96.7b]:       "När du betalar vägtullar, kom ihåg att det är nödvändigt att frigöra        kvartal en full 3 sekunder innan de passerar korgen om du är        reser mer än 60 MPH. "[110,13]:       "När du reser på en enkelriktad gata, stanna till höger, så att inte        störa mötande trafik. "
		-- Leo Kessler

%
Jag antar att en del av variationen mellan Boston förare och resten avland beror på den progressiva Massachusetts förarutbildning Manual somJag råkar ha i min topp skrivbordslåda. Några av de tips för bättre körningär värt att överväga, nämligen:[173.15b]:"När konkurrensen om en vägsträcka eller en parkeringsplats, kom ihåg        att fordonet är i behov av de mest karosseri har rätt-of-way. "[141.2a]:       "Även om det är helt och hållet möjligt att montera en 6 'bil in i en 6'        parkeringsplats, är det sällan möjligt att montera en 6 "bil i        5 'parkeringsplats. "[105,31]:       "Teenage förare tror att de är odödliga, och kör därefter.        Dock bör du undvika frestelsen att bevisa att de har fel. "
		-- Leo Kessler

%
Jag värdesätter vänlighet mot människor först och främst, och vänlighet mot djur. jaginte respekterar lagen, Jag har en total respektlöshet för något anslutnamed samhället utom det som gör vägarna säkrare, öl starkare,maten billigare, och gamla män och kvinnor varmare på vintern, och lyckligarepå sommaren.
		-- Brendan Behan

%
Idaho statens lag gör det olagligt för en man att ge sin kärestaen låda med godis som väger mindre än femtio pounds.
		-- Brendan Behan

%
Om en jury i en rättegång håller utkik efter mer än tjugofyra timmar, detär säker på att rösta frikännande, utom i de fall där det röstar skyldig.
		-- Joseph C. Goulden

%
Om en man hålla sig borta från sin fru för sju år, förutsätter lagen attseparation ha dödat honom; men enligt vår dagliga erfarenhet,det kan mycket väl förlänga sitt liv.
		-- Charles Darling, "Scintillae Juris", 1877

%
"Om en gång en man skämmer sig i mord, mycket snart kommer han att tänkalite av råna; och från råna han nästa kommer att dricka ochSabbats bryta, och från den till ohövlighet och förhalning. "
		-- Thomas De Quincey (1785 - 1859)

%
Om reportrarna inte vet att sanningen är plural, de borde vara advokater.
		-- Tom Wicker

%
Om det fanns en skola för, säg, plåtslagare, som efter treår kvar sina studenter som oförberedda för sina karriärer som gör lagskola, skulle läggas ned i en minut, och utan tvekan av advokater.
		-- Michael Levin, "The Socratic Method"

%
I "Kung Henrik VI, del II," Shakespeare har Dick Butcher föreslåhans kolleger anti-establishment packet-rousers, "Det första vi gör, låt ossdöda alla advokater. "Det åtgärd kan vara extrema, men en liknande känslauttrycktes av Thomas K. Connellan, ordförande för ledningsgruppen, Inc.Tala med företagsledare i Chicago och citerade i Automotive News,Connellan tillskrivas ett mått på USA: s fallande produktivitet till ett överskottav advokater och revisorer, samt en brist på produktion experter. advokateroch revisorer "inte göra det ekonomiska cirkel något större, de bara siffrahur kakan blir uppdelad. Varken yrke ger något mervärdetill produkt. "Enligt Connellan har högproduktiv japanska samhället10 jurister och 30 revisorer per 100.000 invånare. USA har 200advokater och 700 revisorer. Detta tyder på att "den amerikanska andelenPie-bagare och paj-delare är vägen ut ur whack. "Kunde Dick Butcher harvarit en effektivitetsexpert?
		-- Motor Trend, May 1983

%
I Blythe, Kalifornien, förklarar en stad förordning att en person måste ägaåtminstone två kor innan han kan bära cowboystövlar offentligt.
		-- Motor Trend, May 1983

%
I Boston, är det olagligt att hålla groda Jump tävlingar på nattklubbar.
		-- Motor Trend, May 1983

%
I Columbia, Pennsylvania, är det mot lagen för en pilot att kittlaen kvinnlig flygande studenten under hakan med en dammvippa föratt få hennes uppmärksamhet.
		-- Motor Trend, May 1983

%
I Corning, Iowa, det är en förseelse för en man att be sin fru att ridai motorfordon.
		-- Motor Trend, May 1983

%
I Denver är det olagligt att låna din dammsugare till din granne.
		-- Motor Trend, May 1983

%
I Devon, Connecticut, är det olagligt att gå baklänges efter solnedgången.
		-- Motor Trend, May 1983

%
I Greene, New York, är det olagligt att äta jordnötter och gå bakåt påtrottoarer när en konsert är på.
		-- Motor Trend, May 1983

%
I Lexington, Kentucky, är det olagligt att bära en glasstrut i fickan.
		-- Motor Trend, May 1983

%
I Lowes Crossroads, Delaware, är det ett brott mot lokal lagstiftning för varjepilot eller passagerare att bära en glasstrut i fickan medanantingen flyga eller väntar på att gå ombord på ett plan.
		-- Motor Trend, May 1983

%
I Memphis, Tennessee, är det olagligt för en kvinna att köra en bil omDet är en man antingen kör eller går framför det vifta med en rödflagga för att varna närmar bilister och fotgängare.
		-- Motor Trend, May 1983

%
I Ohio, om du ignorerar en talare på dekoration dag till en sådan omfattningatt offentligt spela krocket eller beckhäst inom en mil avtalarens monter, kan du dömas till böter $ 25.00.
		-- Motor Trend, May 1983

%
I Pocataligo, Georgien, är det ett brott för en kvinna över 200 poundsoch klädd i shorts pilot eller rida i ett flygplan.
		-- Motor Trend, May 1983

%
I Pocatello, Idaho, en lag som antogs 1912 under förutsättning att "Det redovisadedolda vapen är förbjudet, om inte samma ställs ut till allmänheten. "
		-- Motor Trend, May 1983

%
I Seattle, Washington, är det olagligt att bära ett dolt vapen somär över sex fot i längd.
		-- Motor Trend, May 1983

%
I Tennessee är det olagligt att skjuta något annat spel än valar från enrörliga bil.
		-- Motor Trend, May 1983

%
Förr i världen i England, kan du vara hängd för att stjäla ett får eller enbrödlimpa. Men om ett får stal en limpa bröd och gav den tilldig, skulle du endast prövas för mottagning, ett brott belagt med fyrtiofransar med katten eller hunden, beroende på vilket som var praktiskt. Om du stal en hundoch fångades, du straffas med tolv kanin slag, även om detvar svårt att hitta kaniner tillräckligt stora eller tillräckligt starka för att slå dig.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
I Tulsa, Oklahoma, är det mot lagen att öppna en läsk flaska utanöverinseende av en licensierad ingenjör.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
I West Union, Ohio, kan Ingen gift man gå flyga utan sin maketillsammans när som helst, om han har varit gift i mer än 12 månader.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Det har länge varit märkt att juryer är skoningslösa för rån och full avseende för barnamord. En intressant fråga, min kära Sir! jurynär rädd för att bli rånad och har passerat den ålder då det kan vara ett offerav barnamord.
		-- Edmond About

%
Det är mot lagen för ett monster för att ange gränserna för företagensUrbana, Illinois.
		-- Edmond About

%
Det är olagligt att köra ner mer än två tusen får HollywoodBoulevard på en gång.
		-- Edmond About

%
Det är olagligt att säga "Åh, Boy" i Jonesboro, Georgien.
		-- Edmond About

%
Det är Mr Mellon credo som $ 200.000.000 kan göra något fel. Vårbrott består i att ifrågasätta den.
		-- Justice Robert H. Jackson

%
Det är Texas lag som när två tåg möter varandra vid en järnvägsövergång,varje ska komma till en punkt, och ingen skall fortsätta tills den andrahar gått.
		-- Justice Robert H. Jackson

%
Det verkar dessa två killar, George och Harry, som anges i en Hot Airballong för att korsa USA. Efter fyrtio timmar i luften, Georgevände sig till Harry, och sa, "Harry, jag tror att vi har kommit ur kurs! Vimåste ta reda på var vi är. "Harry kyler luften i ballongen, och de stiger ned till undermolntäcke. Långsamt glider över landskapet, fläckar George en manstår under dem och skriker ut, "Ursäkta mig! Kan du berättadär vi är?"Mannen på marken skriker tillbaka, "Du är i en ballong, ungefärfemtio fot i luften! "George vänder sig till Harry och säger: "Ja, det man * måste * vara en advokat".Svar Harry, "Hur kan du säga?"."Eftersom den information han gav oss är 100% korrekt, och totaltonyttig!"Det är slutet av skämtet, men för er som fortfarande är oroligGeorge och Harry: de hamnar i drycken, och göra framsidan avNew York Times: "Balloonists dränkts av advokat".
		-- Justice Robert H. Jackson

%
Det ska vara olagligt för någon misstänkt person att vara inom kommunen.
		-- Local ordinance, Euclid Ohio

%
Det är olagligt i Wilbur, Washington, att rida en ful häst.
		-- Local ordinance, Euclid Ohio

%
Det nyligen kommit till Fortune uppmärksamhet som forskarna har slutatanvändning av laboratorieråttor till förmån för advokater. Verkar som det finns intebara mer av dem, men du inte får så känslomässigt fäst. Det endasvårighet är att det ibland är svårt att tillämpa det experimentellaresultat för människor.[Det finns också vissa saker även en råtta inte kommer att göra. Ed.]
		-- Local ordinance, Euclid Ohio

%
Domare, som klass, display, i fråga om att arrangera underhållsbidrag, attvårdslös generositet som finns endast hos män som ger bortnågon annans pengar.
		-- P. G. Wodehouse, "Louder and Funnier"

%
Kom bara ihåg: när du går till domstol, du lita på ditt öde tilltolv personer som inte var smart nog att komma ut ur juryarbetsuppgift!
		-- P. G. Wodehouse, "Louder and Funnier"

%
Kansas State lagen kräver fotgängare korsar vägar på natten för attbära bakljus.
		-- P. G. Wodehouse, "Louder and Funnier"

%
Kirkland, Illinois, förbjuder lag bin att flyga över byn eller genomnågon av dess gator.
		-- P. G. Wodehouse, "Louder and Funnier"

%
Vet hur man sparar 5 drunknings advokater?-- Nej?BRA!
		-- P. G. Wodehouse, "Louder and Funnier"

%
Lagar är som korv. Det är bättre att inte se dem som görs.
		-- Otto von Bismarck

%
Lagstiftningen föreslås i Illinois delstatsparlament, maj 1907:"Speed ​​på länsvägar kommer att begränsas till tio miles i timmenom bilisten ser en fogde som inte verkar ha haft endricka i 30 dagar, när föraren kommer att tillåtas att göra vad han kan. "
		-- Otto von Bismarck

%
Låt oss komma ihåg att vår är en nation av advokater och ordning.
		-- Otto von Bismarck

%
Låt oss säga att din vigselring faller i brödrosten, och när du hållerhanden för att hämta det, du lider smärta och lidande samtPsykiskt lidande. Du skulle stämma:* Brödrost tillverkare, för underlåtenhet att i instruktionerna  avsnitt som säger att du ska aldrig aldrig aldrig någonsin hålla dig hand  i brödrosten, påståendet "Inte ens om din vigselring faller  där inne".* Butiken där du köpte brödrost, för att sälja den till ett självklart  cretin som själv.* Union Carbide Corporation, vilket inte är direkt ansvarig i detta  fallet, men som känner så skyldig att det förmodligen skulle skicka dig  en stor kontantavräkning ändå.
		-- Dave Barry

%
... Logiskt osammanhängande, semantiskt obegriplig, och lagligt ...oklanderlig!
		-- Dave Barry

%
Loud rapningar när hon gick runt flygplatsen är förbjudet i Halstead, Kansas.
		-- Dave Barry

%
Marijuana är lagligt en dag, eftersom många juridikstudentersom nu röker hasch dag kommer att bli kongress och legaliseradet för att skydda sig själva.
		-- Lenny Bruce

%
Män tror ofta - eller låtsas - att "lagen" är något heligt, elleråtminstone en vetenskap - en ogrundad antagande mycket bekvämt att regeringar.
		-- Lenny Bruce

%
Minderåriga i Kansas City, Missouri, är inte tillåtet att köpa knallpulverpistoler;de kan köpa hagelgevär fritt, dock.
		-- Lenny Bruce

%
Aldrig skjuta upp till i morgon vad du kan göra idag. Det kan finnas enlag mot det vid denna tidpunkt.
		-- Lenny Bruce

%
ALDRIG väja att träffa en advokat cykla - det kan vara din cykel.
		-- Lenny Bruce

%
New Hampshire lag förbjuder dig att utnyttja dina fötter, nicka, eller inågot sätt hålla takt med musiken i en krog, restaurang eller café.
		-- Lenny Bruce

%
Av ______ Naturligtvis är det mordvapnet. Vem skulle rama in någon med en falsk?
		-- Lenny Bruce

%
Gamla Barlow var en korsning betalningsmedel vid en korsning där ett expresstågrevs en bil och dess passagerare. Att vara huvudvittne, hansvittnesmål var oerhört viktigt. Barlow förklarade att natten var mörkt,och han viftade lykta frenetiskt, men föraren av bilen betalatsingen uppmärksamhet till signalen.Järnvägföretaget vann målet, och VD för företagetkompletterat gamling för hans berättelse. "Du gjorde underbart", sade han,"Jag var rädd att du skulle tveka i vittnesbörd.""No sir", utropade äldre ", men jag var säker rädd att durnedadvokat tänkte fråga mig om min lykta tändes "
		-- Lenny Bruce

%
När han hade ena benet i Vita huset och nationen darrade under hansbrusar. Nu är han en SKRUTTIG påve i Coca-Cola bälte och en bror tillgivna pastorer som belabor halfwits i galvaniserat järn hyddor bakomjärnvägen varven. "ombud för supportrar av Tennessee anti-evolutionlag på omfattningar "Monkey Trial" i 1925.
		-- H. L. Mencken, writing of William Jennings Bryan,

%
... Vår andra helt sant nyhet skickades till mig av Mr H. BoyceConnell Jr i Atlanta, Ga., Där han är inblandad i en advokatbyrå. En sakJag tycker om South är folk där bryr sig om tradition. Om någonblir överlämnade ett namn som "H. Boyce," han hänger på det, lägger det på sin juridiskabrevpapper, även skickar den till sin son, snarare än att göra vad en mindre människaskulle göra, såsom få det ändrat eller döda sig själv.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh förarens test(10) Potholes är(A) extremt farlig.(B) patriotisk.(C) fel av den tidigare administrationen.(D) alla kommer att fastställas nästa sommar.Rätt svar är (b). Potthål förstöra opatriotiskt, unamerican,importerade bilar, eftersom hålen är större än bilarna. Om du kör enstor, patriotisk, amerikansk bil du har inget att oroa sig för.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh förarens test(2) Ett trafikljus vid en korsning ändras från gult till rött, bör du(A) sluta omedelbart.(B) gå långsamt genom korsningen.(C) blåsa hornet.(D) golvet.Rätt svar är (d). Om du sa (c), du var nästan rätt, såge dig själv en halv punkt.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh förarens test(3) När du stannar vid en korsning bör du(A) se trafikljuset för ditt körfält.(B) titta på fotgängare korsar gatan.(C) blåsa hornet.(D) se trafikljus för den korsande gatan.Rätt svar är (d). Du måste börja så snart trafikljusetför den korsande gatan blir gul. Svar (c) är värt en halv punkt.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh förarens test(4) Avgas är(A) välgörande.(B) inte skadligt.(C) giftiga.(D) ett punkband.Rätt svar är (b). Den inblandning Washington eco-freak kommunistbyråkrater som säger något annat ljuger. (Meddelande till dem som svarade (d).Gå tillbaka till Kalifornien där du kom ifrån. Din slag är inte välkomna här.)
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh förarens test(5) Din bil horn är en viktig del av säkerhetsutrustning. Hur ofta bördu testa det?(A) en gång om året.(B) en gång i månaden.(C) en gång dagligen.(D) en gång i timmen.Rätt svar är (d). Du bör testa bilens horn åtminstone en gångvarje timme, och oftare på natten eller i bostadsområden.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh Förar Test(7) Bilen direkt framför dig har en blinkande rätt baklykta    men en stadig vänster baklykta. Det betyder(A) en av bakljus är bruten; du ska blåsa ditt hornatt ringa problemet till förarens uppmärksamhet.(B) föraren signalerar en högersväng.(C) föraren signalerar en vänstersväng.(D) föraren ut ur staden.Rätt svar är (d). Bakljus används i vissa utländskaländer för att signalera svängar.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh Förar Test(8) Fotgängare är(A) irrelevant.(b) kommunister.(C) en olägenhet.(D) svårt att rensa bort frontgallret.Rätt svar är (a). Fotgängare är inte i bilar, så de ärhelt irrelevant för körning; du ska ignorera dem helt.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Pittsburgh förarens test(9) Vägar saltas för att(A) döda gräs.(B) smälta snö.(C) hjälpa ekonomin.(D) förhindra gropar.Rätt svar är (c). Väg saltning sysselsätter tusentals personerdirekt, och miljontals mer indirekt, exempelvis salt gruvarbetare ochrustproofers. Viktigast minskar saltning livslängden för bilar,och därmed främja bil- och stålindustrin.
		-- Dave Barry, "This Column is Nothing but the Truth!"

%
Hon grät, och domaren torkade tårarna med min checkhäfte.
		-- Tommy Manville

%
Sho "de måste ha det mot lagen. Skjuta, ever'body git hög,de skulle inte finnas någon git upp och mata kycklingarna. Hihi.
		-- Terry Southern

%
Vissa män är heterosexuella, och vissa är bisexuella och vissa män tror inteom sex alls ... de blir advokater.
		-- Woody Allen

%
Några av de mest intressanta dokument från Sveriges medeltid ärgamla läns lagar (bra, vi aldrig haft länen men det är närmast motsvarandeJag kan hitta för "Landskap"). Dessa lagar har skrivits ned någon gång i13-talet, men går tillbaka ända ned till vikingatiden. Den äldsta ärvästgöta lag som tydligt har hedniska influenser, tunt täckt med någonChristian stuff. I denna lag, finner vi en sida om "Lekare", som är denFornnordiska ordet för en artist, skådespelare / gycklare / musiker etc. Här ären automatisk översättning, där jag har skrivit "artist" som motsvarar"Lekare"."Om en konstnär är slagen, ska ingen betala böter för det. Om en konstnärär skadade, en sådan som går med hurdie-gurdie eller reser medfiol eller trumma, då människor ska ta en vild kviga och föraut på en sluttning. Då skall de raka bort allt hår frånkviga svans, och smörj svansen. Sedan konstnären skall gesnyligen smord skor. Sedan skall han ta tag i kviga svans,och en man ska slå den med en skarp piska. Om han kan hålla henne, hanskall ha djuret. Om han inte kan hålla henne, skall han uthärda vadhan fick, skam och sår. "
		-- Woody Allen

%
Ibland kan en man som förtjänar att ses ned på grund av att han är endåre föraktas bara för att han är en advokat.
		-- Montesquieu

%
Texas lag förbjuder någon att ha en tång i sin ägo.
		-- Montesquieu

%
Djuren är inte så dum som man tror - de har varkenläkare eller advokater.
		-- L. Docquier

%
Arkansas lagstiftaren antagit en lag som säger att ArkansasRiver kan stiga högre än till Main Street bron i Little Rock.
		-- L. Docquier

%
Staden Palo Alto, i sin officiella beskrivningen av parkeringsplats standarder,anger graden av rullstols ramper i termer av centimeterstiga per fot körning. En kompromiss, jag kan tänka mig ...
		-- L. Docquier

%
Skillnaden mellan en advokat och en tupp är atttupp stiger upp på morgonen och clucks trots.
		-- L. Docquier

%
District of Columbia har en lag som förbjuder dig att utöva påtryckningar påen ballong och därigenom orsaka ett visslande ljud på gatorna.
		-- L. Docquier

%
Domaren ålade jaywalker femtio dollar och berättade för honom om han varfångas igen, skulle han kastas i fängelse. Fin idag, svalare i morgon.
		-- L. Docquier

%
Motiveringarna till drogtester är en del av den för närvarande fashionabladebatt om att återställa USA: s "konkurrenskraft." Läkemedel, har det varitavslöjat, är ansvariga för skenande frånvaro, minskad produktion och dåligkvalitetsarbete. Men är drogtestning i själva verket på ett rationellt sätt i samband meduppståndelse konkurrenskraft? Kommer laddning atmosfären iarbetsplats med rädslan för utsöndrings svek ärligt sporra produktivitet?Mycket buller har gjorts om rehabilitering arbetaren använda droger, menhittills de allra flesta program avslutas med enkel bränning eller inteuthyrning av förövaren. Denna praxis kan förvärra, inte lindra dennationens produktivitetsproblem. Om den ekonomiska rehabiliteringen är den ultimataMålet med drogtestning, då kriterier överge rehabilitering avnarkotikaanvändande arbetare är den renaste av hyckleri och det värsta av rationalisering.Fjärde rättelse och drogtestning på arbetsplatsen, "Tim Moore, Harvard Journal of Law & Public Policy, vol.10, nr 3 (sommar 1987), sid. 762-768.
		-- The concluding paragraph of "Constitutional Law: The

%
Lagen, i sin majestätiska jämlikhet, förbjuder de rika, liksom de fattiga,att sova under broarna, att tigga på gatorna, och att stjäla bröd.
		-- Anatole France

%
Den lagstiftare, av alla varelser, beror de flesta lagen trohet. Han av alla mänbör bete sig som om lagen tvingade honom. Men det är den universellasvaghet för mänskligheten att det vi får till administrera vi nu föreställavi äger.
		-- H. G. Wells

%
Den minst framgångsrika Equal Pay Annons1976 pekade Europeiska ekonomiska gemenskapen ut till den irländskaRegeringen att det ännu inte hade genomfört de överenskomna jämställdhet mellan könenlagstiftning. Dublin regeringen omedelbart annonseras för en lika lönkronofogden. Annonsen erbjuds olika löneskalor förmän och kvinnor.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Straffet för skratt i en rättssal är sex månader i fängelse; om detinte för detta straff, juryn skulle aldrig höra bevis.
		-- H. L. Mencken

%
De befogenheter inte delegeras till Förenta staterna av konstitutionen, ellerförbjudet enligt den till stater, reserveras till stater respektive,eller till folket.
		-- U.S. Constitution, Amendment 10. (Bill of Rights)

%
Den primära förutsättning för varje ny skattelagstiftning är att det ska undanta tillräckligtväljarna att vinna nästa val.
		-- U.S. Constitution, Amendment 10. (Bill of Rights)

%
Staten lag Pennsylvania förbjuder sjunga i badkaret.
		-- U.S. Constitution, Amendment 10. (Bill of Rights)

%
Värsta JuryEn mordrättegång i Manitoba i februari 1978 var långt, nären jurymedlem avslöjade att han var helt döv och inte haravlägsna aning om vad som hände.Domaren, Mr Justice Solomon, frågade honom om han hade hört någonbevis alls och, när det inte fanns något svar, avskedade honom.Spänningen som detta orsakade endast motsvarade när en andrajurymedlem avslöjade att han talade inte ett ord engelska. En flytande franskahögtalare, uppvisade han stor överraskad när berättade, efter två dagar, att hanhörde en mordrättegång.Försöket övergavs när en tredje jurymedlem sade att han ledfrån båda villkor, samtidigt som OBEVANDRAD på engelskaoch nästan lika döv som den första jurymedlem.Domaren beordrade en ny rättegång.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Det finns en Massachusetts lag som innebär att alla hundar har bakbenenbundet under april månad.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Det finns inget bättre sätt att utöva fantasin än studiet av lagen.Ingen poet som har tolkat naturen så fritt som en jurist tolkar sanningen.
		-- Jean Giraudoux, "Tiger at the Gates"

%
Det råder ingen tvekan om att min advokat är ärlig. Till exempel, när hansparade hans självdeklaration förra året, förklarade han halva sin lönsom "kapitalinkomst."
		-- Michael Lara

%
"Det var en intressant utveckling i CBS-Westmoreland rättegången:båda sidor överens om att efter rättegången skulle Andy Rooney tillåtasprata med juryn för tre minuter om små saker som irriterade honomunder rättegången. "
		-- David Letterman

%
Det finns ingen rättvisa i världen.New York åklagare Thomas Dewey efter Luciano hadesparade Dewey från mordet av den holländska Schultz (genom att beställamordet på Schultz istället)
		-- Frank Costello, on the prosecution of "Lucky" Luciano by

%
Virginia lag förbjuder badkar i huset; baljor måste hållas på gården.
		-- Frank Costello, on the prosecution of "Lucky" Luciano by

%
Vi kanske inte gillar läkare, men åtminstone de läkare. Bankers är aldrigpopulär men åtminstone de bank. Policeman polisen och begravnings taunder. Men advokater inte ge oss rätt. Vi får inte glädjerik ljusi rättsvetenskap, utan prejudikat, invändningar, överklaganden, stag,anmälningar och blanketter, motioner och kontra rörelser, alla på $ 250 en timme.
		-- Nolo News, summer 1989

%
Vi måste inse att en stad är bättre med dåliga lagar, så länge deförblir fast, sedan med bra lagar som ständigt förändras, attavsaknaden av lärande i kombination med ljud sunt förnuft är mer användbar änden typ av skicklighet som spårar ur, och att som en allmän regel,stater bättre styrs av mannen på gatan än av intellektuella.Dessa är den typ av människor som vill synas klokare än de lagar somvill få sin egen väg i varje allmän diskussion, eftersom de anser attde kan inte visa upp sin intelligens i fråga om större betydelse, ochsom följd, mycket ofta ta ruin på deras land.
		-- Cleon, Thucydides, III, 37 translation by Rex Warner

%
Välkommen till Utah.Om du tror att våra sprit lagar är roligt, bör du se vår underkläder!
		-- Cleon, Thucydides, III, 37 translation by Rex Warner

%
Vad har du när du har sex advokater begravd upp till halsen i sanden?Inte nog sand.
		-- Cleon, Thucydides, III, 37 translation by Rex Warner

%
När varnas för ett intrång av pinglande glas eller på annat sätt, en) Lugnsjälv 2) Identifiera inkräktaren 3) Om fientlig, döda honom.Steg nummer tre är av särskild betydelse. Om du lämnar killen levandeav missriktad softheartedness, kommer han att betala din generositetgenom att stämma dig för att ha orsakat hans efterföljande paraplegi och försöka tvinga digför att stödja honom för resten av sitt ruttna liv. I domstol han åberopaatt han var deprimerad eftersom samhället hade svikit honom, och att han varsöker Moder Teresa för komfort och att erbjuda sina tjänster tillfattig. I rättegången, kommer du att förlora. Om, å andra sidan, du dödarhonom, är det mesta som du kan förvänta sig att en släkting kommer att medföra en felaktigdöd åtgärder. Du kommer att ha två fördelar: för det första, bara det finnas dinberättelse; glömma Moder Teresa. För det andra, även om du förlorar, hur mycket skullebum liv vara värt ändå? Mycket mindre än 50 år till ett värde avförlamning. Inte spela George Bush och Saddam Hussein. Avsluta jobbet.
		-- G. Gordon Liddy's "Forbes" column on personal security

%
Om det är en plikt att dyrka solen är ganska säker på att vara ett brott attgranska lagar värme.
		-- Christopher Morley

%
Varför en likbil häst snicker, dragande en advokat bort?
		-- Carl Sandburg

%
Varför New Jersey har mer giftiga avfallsdeponier och Kalifornien harfler advokater?New Jersey hade förstahandsval.
		-- Carl Sandburg

%
Med kongressen, varje gång de gör ett skämt det är en lag; och varje gångde gör en lag det är ett skämt.
		-- Will Rogers

%
"Visst, om en enskild stoppades och anklagades för snatteri efter promenader i Neiman-Marcus de förväntar sig att bli så småningom berättade vad de stal allegedly. Det vore absurt om en officer att berätta den tilltalade att "du vet vad du stal jag inte berätta." Eller att helt enkelt lämna den anklagade en katalog över Neiman-Marcus hela inventering och säga "det är där någonstans, räkna du ut det." "    - Domaren Brooke Wells att fatta i del IBMs Motion för att begränsa       SCO: s krav
		-- Will Rogers

%
"Obligatorisk enande yttrande uppnår endast genom enhälligt beslut av kyrkogård."    - Rättvisa Jackson, skriva för de flesta, i West Virginia       State Board of Education v. Barnette 319 US 624 nr 591
		-- Will Rogers

%
"Om det finns någon fixstjärna i vår konstitutionella konstellation, är det att ingen officiell, hög eller ringa, kan ordinera vad som skall ske ortodox i politik, nationalism, religion, eller andra frågor av åsikt eller tvinga medborgarna att erkänna med ord eller handla sin tro däri. Om det finns några omständigheter som medger ett undantag, de inte nu inträffa till oss."    - Rättvisa Jackson, skriva för de flesta, i West Virginia       State Board of Education v. Barnette 319 US 624 nr 591
		-- Will Rogers

%
"Rätten till tanke- och religionsfrihet som garanteras av Konstitution mot statliga åtgärder omfattar både rätten att tala fritt och rätten att avstå från att tala alls, utom i den mån som viktiga operationer regerings kan kräva det för bevarandet av en ordnad samhälle --- som i fallet med tvång till vittna i domstol. "    - Rättvisa Murphy, i concurrance, West Virginia State Board of       Utbildning v. Barnette 319 US 624 nr 591
		-- Will Rogers

%
