  Lite smärta aldrig skadat någon.
		-- Arthur Baer, American comic and columnist

%
  "En enhetlig, neutral Tyskland? Med tanke på att nationens kulturarv, en sådan  fras kan visa sig vara oxymoron av decenniet. "-Kevin M.  Matarese, Fulda, Västtyskland; såsom framgår av "Letters", Tid  tidskrift, s. 5 den 5 mars 1990.
		-- Arthur Baer, American comic and columnist

%
  Ett muntligt avtal är inte värt papperet det är skrivet på. Omfatta  mig. -Samuel Goldwyn
		-- Arthur Baer, American comic and columnist

%
  Kristus föddes 4 f.Kr.
		-- Arthur Baer, American comic and columnist

%
  Cum tacent, LARMANDE. När de är tysta, de skriker. -Cicero
		-- Arthur Baer, American comic and columnist

%
  Mina herrar, jag vill att du ska veta att jag inte alltid rätt, men jag är  aldrig fel. -Samuel Goldwyn
		-- Arthur Baer, American comic and columnist

%
  Goes (Gick) över som en ledande ballong.
		-- Arthur Baer, American comic and columnist

%
  Tuta, om du är emot buller!
		-- Arthur Baer, American comic and columnist

%
  Jag ska ge dig en bestämd kanske. -Samuel Goldwyn
		-- Arthur Baer, American comic and columnist

%
  Jag tänker inte säga, "jag sa."
		-- Arthur Baer, American comic and columnist

%
  Jag är en djupt ytlig person. -Andy Warhol
		-- Arthur Baer, American comic and columnist

%
  Jag är stolt över min ödmjukhet.
		-- Arthur Baer, American comic and columnist

%
  Jag kan motstå allt utom frestelser. -Oscar Wilde
		-- Arthur Baer, American comic and columnist

%
  Om Roosevelt levde, skulle han vända sig i sin grav. -Samuel  Goldwyn
		-- Arthur Baer, American comic and columnist

%
  Om jag kunde släppa död just nu, skulle jag vara den lyckligaste mannen vid liv!
		-- Samuel Goldwyn

%
  Om du faller och bryter benen, inte komma springande till mig. -Samuel  Goldwyn
		-- Samuel Goldwyn

%
  Jag har aldrig sätta på sig ett par skor tills jag har burit dem fem år.
		-- Samuel Goldwyn

%
  Det är inte en optisk illusion. Det ser ut precis som en.
		-- Samuel Goldwyn

%
  Det är mer än magnifik, det är mediokra. -Samuel Goldwyn
		-- Samuel Goldwyn

%
  Får jag ställa en fråga?
		-- Samuel Goldwyn

%
  Ingen går till den restaurangen längre, det är alltid alltför trångt.  (Skrivs Yogi Berra)
		-- Samuel Goldwyn

%
  Våra komedier är att inte bli utskrattad. -Samuel Goldwyn
		-- Samuel Goldwyn

%
  Avstickning är sådan söt sorg. -William Shakespeare
		-- Samuel Goldwyn

%
  Förhalning innebär aldrig behöva säga att du är ledsen.
		-- Samuel Goldwyn

%
  "Professionell certifiering för bil människor kan låta som en  oxymoron. "-The Wall Street Journal, sida B1, tisdag den 17 juli  1990.
		-- Samuel Goldwyn

%
  Med hänvisning till en bok: Jag läste en del av det hela vägen igenom.
		-- Samuel Goldwyn

%
  Rökning är den vanligaste orsaken till statistiken.
		-- Samuel Goldwyn

%
  Vissa ungkarlar vill ha en meningsfull över natten förhållande.
		-- Samuel Goldwyn

%
  Att tala om en bit av film dialog: Låt oss ha några nya  klichéer. -Samuel Goldwyn
		-- Samuel Goldwyn

%
  Scenen är tråkig. Säg till honom att lägga mer liv i sin döende.
		-- Samuel Goldwyn

%
  Tack och lov Jag är ateist.
		-- Samuel Goldwyn

%
  Denna rapport är fylld med brister.
		-- Samuel Goldwyn

%
  Vi är inte att föregripa eventuella nödsituationer.
		-- Samuel Goldwyn

%
  Vi utbetala honom, men han är värd det. -Samuel Goldwyn
		-- Samuel Goldwyn

%
  Hans ära rotad i vanära stod  Och tro otrogen höll honom falskt sant.
		-- Alfred Lord Tennyson

%
  Den goda oxymoron, för att definiera den genom en själv illustration, måste vara en  planerade OVARSAMHET. -Wilson Follett
		-- Alfred Lord Tennyson

%
  En irländare är aldrig i fred utom när han kämpar.
		-- Alfred Lord Tennyson

%
  Jag förundras över styrkan i mänsklig svaghet.
		-- Alfred Lord Tennyson

%
  Alltid vara ärlig, även när du inte menar det. -Irene Peter
		-- Alfred Lord Tennyson

%
  Leva inom din inkomst, även om du måste låna för att göra det.
		-- Josh Billings

%
  Naturligtvis kan jag hålla hemligheter. Det är människorna jag berätta för dem att det  kan inte hålla dem. -Anthony Haden-Guest
		-- Josh Billings

%
  Det bästa botemedlet mot sömnlöshet är att få mycket sömn. -W. C. Fält
		-- Josh Billings

%
  Jag minns tydligt att glömma det. -Clara Barton
		-- Josh Billings

%
  Vi måste tro på fri vilja. Vi har inget annat val. -Isaac B. Singer
		-- Josh Billings

%
  Jag skulle ge min högra arm att vara ambidextrous.
		-- Josh Billings

%
  Monoteism är en gåva från gudarna.
		-- Josh Billings

%
  Efter att de blev av med dödsstraff, var de tvungna att hänga två gånger  så många människor som tidigare.
		-- Josh Billings

%
  Jag har aldrig gillat dig, och jag kommer alltid. -Samuel Goldwyn
		-- Josh Billings

%
  Varför inte koppla `em up i treor? -Yogi Berra
		-- Josh Billings

%
  Våra likheter är olika. -Dale Berra, son till Yogi
		-- Josh Billings

%
  Efter Donald Trumps stretch limousine stals och hittades  oskadad några kvarter bort; sade han, "Ingenting var stulet. Jag hade  en ärlig tjuv "-. International Herald Tribune, sidan 3, den 2 mars  1992
		-- Josh Billings

%
  Vissa fågelpopulationer skyhöga ner-Headline Av en artikel iScience News, sid 126, 20 februari, 1993.
		-- Josh Billings

%
  De flesta bakterier ha anständigheten att vara mikroskopisk. Epulopiscium  fishelsoni är inte bland dem. Den nyligen identifierade en encelliga  makromikroorganismen är en full .5 mm lång, tillräckligt stora för att ses  med blotta ögat. Beskrivs i den aktuella Nature, "Det är en  miljoner gånger så stora som en typisk bakterie. "- Time, sidan 25,  29 Mars 1993
		-- Josh Billings

%
  "Triumph utan seger, oredovisade historia persiska  Gulfkriget ", -Headline publicerades i USA News & World Report,  1992.
		-- Josh Billings

%
  En tom hytt drev upp och Sarah Bernhardt kom ut. -Arthur Baer,  Amerikansk komiker och kolumnist
		-- Josh Billings

%
  Hon brukade diet på alla typer av mat hon kunde lägga händerna på.
		-- Arthur Baer, American comic and columnist

%
  Det första villkoret för odödlighet är död. -Stanislaw Lec
		-- Arthur Baer, American comic and columnist

%
  Lika känd som den okända soldaten.
		-- Arthur Baer, American comic and columnist

%
  Jag måste följa människor. Är jag inte deras ledare? -Benjamin Disraeli
		-- Arthur Baer, American comic and columnist

%
  Hegel hade rätt när han sade att vi lär oss av historien att människan  kan aldrig lära sig något av historien. -George Bernard Shaw
		-- Arthur Baer, American comic and columnist

%
  William Safire regler för skrivandet som ses i New York Times     Placera inte uttalanden i negativ form.     Och inte börja meningar med en kombination.     Om du läsa ditt arbete, hittar du på rereading att en stor     många upprepningar kan undvikas genom rereading och redigering.     Använd aldrig en lång ord när en diminutiv kommer att göra.     Okvalificerade superlativ är det värsta av allt.     Om ett ord är olämpligt i slutet av en mening, är en länk verb.     Undvik trendiga talesätt som låter flagnande.     Aldrig, aldrig använda repetitiva uppsägningar.     Undvik också obekväma eller påverkas allitteration.     Sist men inte minst, undvika klyscha är som pesten.
		-- Arthur Baer, American comic and columnist

%
  Alla skriver på väggarna utom mig. -Said Att vara graffiti ses i Pompeii
		-- Arthur Baer, American comic and columnist

%
  Jag snubblade över ett hål som stack upp ur marken.
		-- Arthur Baer, American comic and columnist

%
  Jag tror inte att någon ska skriva sin självbiografi förrän efter  de är döda. -Samuel Goldwyn
		-- Arthur Baer, American comic and columnist

%
  Denna sida har avsiktligt lämnats tom.
		-- Arthur Baer, American comic and columnist

%
  Ondskan är inte alla dåliga.
		-- Arthur Baer, American comic and columnist

%
  Jag håller inte med enhällighet.
		-- Arthur Baer, American comic and columnist

%
  "Det är ett steg framåt även om det fanns inga framsteg."  President Hosni Murbarak Egyptens försök att sätta bästa ansiktet  på en nedslående toppmöte mellan president Clinton och  den syriska diktatorn Hafez Assad.
		-- Arthur Baer, American comic and columnist

%
  "Jag undviker alltid profete förväg eftersom det är mycket bättre  att sia efter händelsen redan har ägt rum. "- Winston  Churchill
		-- Arthur Baer, American comic and columnist

%
 Alla sanningar är sanna för en sträcka, inklusive denna. -XA
		-- Arthur Baer, American comic and columnist

%
 Antag en dygd, om du har det inte. -William Shakespeare
		-- Arthur Baer, American comic and columnist

%
 Alla generaliseringar är farliga, inklusive denna.
		-- Arthur Baer, American comic and columnist

%
