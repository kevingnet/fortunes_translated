En svart katt korsar din väg betyder att djuret går någonstans.
		-- Groucho Marx

%
En vän till mig är i Voodoo akupunktur. Du behöver inte gå.Du ska bara gå ner på samma gata och ... Ooohh, det är mycket bättre.
		-- Steven Wright

%
En stor spindel i ett gammalt hus byggt en vacker bana där för att fånga flugor.Varje gång en fluga landade på webben och intrasslad i det spindeln slukadehonom, så att när en annan fluga kom han skulle tro på nätet var en säker ochlugn plats att vila. En dag en ganska intelligent fluga surrade runtöver banan så länge utan belysning som spindeln dök upp och sa,"Kom ner." Men flugan var för smart för honom och sade, "Jag har aldrig tändadär jag inte ser andra flugor och jag kan inte se några andra flugor i ditt hus. "Så han flög iväg tills han kom till en plats där det fanns en stor många andraflugor. Han var på väg att slå sig ner bland dem när ett bi surrade upp och sade,"Vänta, dum, det är flugpapper. Alla dessa flugor fångas." "Var intedum ", sade fly", de dansar. "Så han lugnat ner sig och fastnadetill flugpapperet med alla andra flugor.Moral: Det finns ingen säkerhet i antal, eller i något annat.
		-- James Thurber, "The Fairly Intelligent Fly"

%
Många människor är rädda för höjder. Inte jag. Jag är rädd för bredder.
		-- Steven Wright

%
En MODERN FABLEAisopos fabler och andra traditionella barns berättelser innebär allegorialltför subtil för dagens ungdom. Barn behöver en uppdaterad meddelandemed samtida omständighet och tomt linje, och tillräckligt kort för att passadagens minuters uppmärksam.Troubled AardvarkEn gång i tiden fanns det en aardvark vars enda glädje i livet varkörning från sin förorts bungalow till sitt jobb på ett stort mäklarfirmai hans nya 4x4. Han hatade sin manipulativ chef, hans beräknande ochoetiska medarbetare, hans giriga hustru, och hans LIPANDE, ogiltigabarn. En dag, Aardvark återspeglas på betydelsen av hans liv ochhans karriär och den okontrollerade, katastrofal minskning med sin nation, desspatetisk ursäkt för ledarskap, och den fullständiga ineffektivitet någonpersonlig insats han kunde göra för att ändra status quo. Övervinnas genom envåg av total depression och självtvivel, bestämde han sig för att ta den endatillvägagångssättet som skulle föra honom ökad komfort och lycka: hankörde till köpcentret och köpte importerade hemelektronikvaror.Sensmoralen i historien: Investera i utländska hemelektronik tillverkare.
		-- Tom Annau

%
En pungråtta måste vara sig själv, och vara sig själv att han är ärlig.
		-- Walt Kelly

%
"En makt så stor, det kan endast användas på gott och ont!"
		-- Firesign Theatre, "The Giant Rat of Summatra"

%
Olyckor orsakar historia.Om Sigismund unbuckle hade tagit en promenad i 1426 och träffade Wat Tyler, denBond Revolt skulle aldrig ha hänt och bilen skulle intehar uppfunnits fram 2026, vilket skulle ha inneburit att all oljakunde ha använts för lampor, vilket sparar den elektriska glödlampan ochwhale, och ingen skulle ha fångat Moby Dick eller Billy Budd.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Alla män är dödliga. Sokrates var dödlig. Därför är alla män är Sokrates.
		-- Woody Allen

%
Alla människor i mitt hus är galen. Killen ovanför mig designsyntetiska hårbollar för keramiska katter. försökte Damen över hallen tillråna ett varuhus ... med en prissättning pistol ... Hon sa, "Ge mig allaav pengarna i valvet, eller jag märkning ner allt i butiken. "
		-- Steven Wright

%
Och nu till något helt annat.
		-- Steven Wright

%
Och nu till något helt densamma.
		-- Steven Wright

%
"Är du säker på att du inte är en encyklopedi försäljare?»Nej, frun. Bara en inbrottstjuv, kommer att plundra lägenheten. "
		-- Monty Python

%
Som poeten sa, "Bara Gud kan göra ett träd" - förmodligen eftersom det ärså svårt att räkna ut hur man får barken på.
		-- Woody Allen

%
Being Ymor högra hand var som försiktigt piskades till döds meddoftande bootlaces.
		-- Terry Pratchett, "The Colour of Magic"

%
Bernard Shaw är en utmärkt människa; Han har inte en fiende i världen, ochingen av hans vänner som han heller.
		-- Oscar Wilde

%
"Boy, tar livet en lång tid att leva."
		-- Steven Wright

%
Bozo är Brotherhood of Dragkedjor och övriga. Bozos är människor som bandtillsammans för skojs skull och vinst. De har inga jobb. Vem som helst som går på entur är en Bozo. Varför en Bozo korsa gatan? Eftersom det finns en Bozopå andra sidan. Den kommer från uttrycket Vos otros, det vill säga andra.De är stora, feta, mitt midja. Den arketyp är en irländsk berusadclown med rött hår och näsa, och blek hud. Fields, William Bendix.Alla tenderar att glida mot Bozoness. Det har Oz i den. de menarväl. De är raka ser förutom att de har uppblåsbara skor. Degillar deras bekvämligheter. De bozos har lärt sig att njuta av sin lediga tid,vilket är hela tiden.
		-- Firesign Theatre, "If Bees Lived Inside Your Head"

%
Men jag alltid sköt in den närmaste backen eller i annat fall, i mörkret.Jag menade inget illa; Jag gillade bara explosionerna. Och jag var noga med att aldrigdödar mer än jag kunde äta.
		-- Raoul Duke

%
"Men jag tycker inte om skräppost !!!!"
		-- Raoul Duke

%
"Men jag vill inte gå på vagnen ...""Åh, inte vara en baby!""Men jag känner mig mycket bättre ...""Nej, du är inte ... i ett ögonblick kommer du att stendöd!"
		-- Monty Python, "The Holy Grail"

%
Förbifarts är enheter som tillåter vissa människor att rusa från punkt A tillpunkt B mycket snabbt medan andra människor rusa från punkt B till punkt A mycketsnabb. Människor som lever vid punkt C, varvid en punkt direkt i mellan, ärofta ges undra vad som är så bra med punkt A som så många människorfrån punkt B är så angelägna om att komma dit och vad som är så bra med punkt Batt så många människor från punkt A är så angelägna om att få _____ där. oftaönskar att folk bara en gång för alla skulle fungera var fande ville vara.
		-- Douglas Adams, "The Hitchhiker's Guide to the Galaxy"

%
Komedi, som medicin, var aldrig tänkt att utövas av allmänheten.
		-- Douglas Adams, "The Hitchhiker's Guide to the Galaxy"

%
Döden svarade inte. Han tittade på SPOLD på samma sätt som en hund serpå ett ben, endast i detta fall det var mer eller mindre tvärtom.
		-- Terry Pratchett, "The Colour of Magic"

%
Inred ditt hem. Det ger en illusion av att ditt liv är merintressant än det egentligen är.
		-- C. Schulz

%
Tror du att när de frågade George Washington för ID som hanbara piskade ut en fjärdedel?
		-- Steven Wright

%
"Kom inte tillbaka förrän du har honom", sade Tick-Tock Man tyst,uppriktigt, extremt farligt.De använde hundar. De använde prober. De använde hjärt platt crossoffs.De använde teepers. De använde mutor. De använde stick tites. De brukadeskrämsel. De använde plåga. De använde tortyr. De använde finks.De använde polisen. De använde husrannsakan och beslag. De använde fallaron. Debegagnade förbättrande incitament. De använde fingeravtryck. De användebertillion systemet. De använde list. De använde svek. De använde förräderi.De använde Raoul-Mitgong men han var inte mycket hjälp. De använde tillämpad fysik.De använde tekniker för kriminologi. Och vad fan, fångade de honom.
		-- Harlan Ellison, "Repent, Harlequin, said the Tick-Tock Man"

%
Ta inte livet så allvarligt, son, är det inte SI OCH SÅ permanent.
		-- Walt Kelly

%
Oroa dig inte om världen närmar sig sitt slut i dag. Det är redan i morgoni Australien.
		-- Charles Schulz

%
Tidigt att stiga, tidigt till sängs, gör en människa frisk, rik och död.
		-- Terry Pratchett, "The Light Fantastic"

%
Eternal intighet är bra om du råkar vara klädd för det.
		-- Woody Allen

%
Eternity är en fruktansvärd tanke. Jag menar, där kommer det att sluta?
		-- Tom Stoppard

%
Ända sedan förhistorisk tid, har vise män försökte förstå vad,exakt, få folk att skratta. Det är därför de kallades "vise män". Allaandra förhistoriska människor var ute punktering varandra med spjut, ochvise män var tillbaka i grottan talesätt: "Hur: Vill du ta minfru? Nej Hur: Här är min fru, ta henne just nu. Nej Hurom: Vill du ta något? Min fru är tillgänglig. No. Hurhandla om ..."
		-- Dave Barry, "Why Humor is Funny"

%
Långt ut i okända bakvatten i omoderna änden avWestern Spiral arm av Galaxy ligger en liten unregarded gul solen.Orbiting detta på ett avstånd av cirka nittio-åtta miljoner miles är enytterst obetydlig liten blågrön planet vars apa-härstammar livformer är så otroligt primitiva att de fortfarande tror digitala klockorär en ganska snyggt idé ...
		-- Douglas Adams, "The Hitchhiker's Guide to the Galaxy"

%
Snabbare, snabbare, du lura, du lura!
		-- Bill Cosby

%
Först några ord om verktyg.I grund och botten är ett verktyg ett objekt som gör att du kan dra nytta avfysikens lagar och mekanik på ett sådant sätt att man allvarligt kan skadasjälv. Idag, människor tenderar att ta verktyg för givet. Om du någonsingående längs gatan och du märker några människor som ser särskiltsjälvbelåten, oddsen är att de tar verktyg för givet. Om jag var du,Jag skulle gå rätt upp och smälla dem i ansiktet.
		-- Dave Barry, "The Taming of the Screw"

%
För min födelsedag fick jag en luftfuktare och en de-luftfuktare ... Jag satte dem ii samma rum och låta dem bekämpa det.
		-- Steven Wright

%
Från det ögonblick tog jag din bok ända tills jag lägger ner var jag skakademed skratt. En dag jag tänker läsa den.
		-- Groucho Marx, from "The Book of Insults"

%
Gud är en komisk spela för en publik som är rädda för att skratta.
		-- Groucho Marx, from "The Book of Insults"

%
Han frågade mig om jag visste vilken tid det var - jag sa ja, men inte just nu.
		-- Steven Wright

%
"Här är något att tänka på: Hur kommer du aldrig se en rubrik som`Psychic vinner lotteri"? "
		-- Jay Leno

%
Hej, vad förväntar ni er från en kultur som * enheter * på * ways * och* Parker * på * uppfarter *?
		-- Gallagher

%
Hög Präst: försvarsmateriel Chapter One, vers nio till tjugosju:Bro. Maynard: Och Saint Attila höjt heliga handgranat upp på högsäger: "O Herre, Välsigna oss detta heliga handgranat, och med detkrossa våra fiender till små bitar. "Och Herren gjorde flin, ochfolk gjorde fest på lammen och hermeliner, och orangutanger, ochfrukostflingor, och Lima bean-Överstepräst: Hoppa lite, broder.Bro. Maynard: Och då Herren talade och sade: "För det första skall tagaut den heliga pin. Då skall du räkna till tre. Inte mer inte mindre.* Tre * skall vara numret på räkningen, och numret påRäkning skall vara tre. * Fyra * skall du inte räkna, och inte hellerräkna du två, förutom att du sedan drager till tre. fem är	RÄTT UT. När antalet tre, varvid det tredje numret nås,då lobbest du din heliga handgranat mot din fiende, som befinnerstygg i mina ögon, skall snus det. Amen.All: Amen.
		-- Monty Python, "The Holy Hand Grenade"

%
"Humor är ett läkemedel som det är på modet att missbruk."
		-- William Gilbert

%
Humorister alltid sitta vid bordet barnens.
		-- Woody Allen

%
Jag är en samvetsgrann man, när jag kastar stenar på sjöfåglar jag lämnar ingen tärnaunstoned.
		-- Ogden Nash, "Everybody's Mind to Me a Kingdom Is"

%
Jag får in abstrakt målning. Real abstrakt - ingen borste, ingen duk,Jag tänker bara om det. Jag gick bara till ett konstmuseum där all konstgjordes av barn. Alla målningarna hängde på kylskåp.
		-- Steven Wright

%
Jag är två med naturen.
		-- Woody Allen

%
Jag argumenterar mycket väl. Fråga någon av mina återstående vänner. Jag kan vinna ett argument påvilket ämne som helst, mot någon motståndare. Folk vet detta, och undvika migparter. Ofta som ett tecken på deras stora respekt, att de inte ens bjuda in mig.
		-- Dave Barry

%
"Jag försäkrar er tanken aldrig ens slagit mig, herre.""I själva verket? Sen om jag var du skulle jag stämma mitt ansikte för förtal."
		-- Terry Pratchett, "The Colour of Magic"

%
Jag grundar min mode smak på vad som inte kliar.
		-- Gilda Radner

%
Jag köpte några begagnade färg. Det var i form av ett hus.
		-- Steven Wright

%
Jag kan inte överbetona betydelsen av god grammatik.Vad en lerkruka. Jag kunde lätt överbetona vikten av godgrammatik. Till exempel kan jag säga: "Dålig grammatik är den vanligaste orsakenlångsam, plågsam död i Nordamerika ", eller" Utan god grammatik, denUSA skulle ha förlorat andra världskriget. "
		-- Dave Barry, "An Utterly Absurd Look at Grammar"

%
"Jag har ändrat mina strålkastare häromdagen. Jag satte i stroboskopljus istället! Nunär jag kör på natten, det ser ut som alla andra står still ... "
		-- Steven Wright

%
Jag kunde dansa med dig tills korna kommer hem. Vid närmare eftertanke jag hellredansa med korna tills du kommer hem.
		-- Groucho Marx

%
Jag förtjänar inte detta pris, men jag har artrit och jag förtjänar inte attantingen.
		-- Jack Benny

%
Jag får inte någon respekt.
		-- Jack Benny

%
Jag dödar inte flugor, men jag gillar att bråka med sina sinnen. Jag håller dem ovanglober. De galen och skrika "Whooa, jag * sätt * alltför hög."
		-- Bruce Baum

%
Jag vill inte leva på i mitt arbete, jag vill leva på i min lägenhet.
		-- Woody Allen

%
Jag slutligen gick till ögonläkare. Jag fick kontakter. Jag behöver bara dem tillläsa, så jag fick flip-ups.
		-- Steven Wright

%
"Jag fick in en hiss i arbetet och den här mannen följde efter mig ... Jagdrivit '1' och han bara stod där ... Jag sa "Hej, vart ska du?" hansa, "Phoenix". Så jag sköt Phoenix. Några sekunder senare dörrarnaöppnat, två tumbleweeds blåste ... vi var i centrala Phoenix. jag tittadepå honom och sa "Du vet, du är den typen av kille jag vill hängamed.' Vi satte sig i bilen och körde ut till sin hydda i öknen.Då ringde telefonen. Han sa "du får det." Jag plockade upp och sa"Hallå?" ... Den andra sidan sa "Är detta Steven Wright?" ... Jag sa "ja ..."Killen sa "Hej, jag är Mr Jones, studielån chef från din bank ...Det verkar som du har missat din sista 17 betalningar, och universitetet dudeltog sade att de fick ingen av de $ 17.000 vi lånade dig ... vivill bara veta vad som hände med pengarna? " Jag sa, "Mr. Jones,Jag ska ge det till dig direkt. Jag gav alla pengar till min vän Slick,och med det han byggde kärnvapen ... och jag skulle uppskatta om du aldrigkallade mig igen. "
		-- Steven Wright

%
Jag fick mitt körkort foto taget ur fokus på ändamålet. NuNär jag får dras över polis ser på det (flytta den närmare ochlängre, försöker se det tydligt) ... och säger: "Här, du kan gå."
		-- Steven Wright

%
Jag fick denna pulveriserad vatten - nu vet jag inte vad jag ska lägga till.
		-- Steven Wright

%
Jag tröttnade på att lyssna på inspelningen på telefonen på filmenteater. Så jag köpte albumet. Jag fick sparkas ut ur en teaternhäromdagen för att föra min egen mat i. hävdade jag att koncessionenstå priserna var upprörande. Dessutom hade jag inte haft en grill i enlänge sedan. Jag gick på teater och tecknet sade vuxna $ 5 barn$ 2,50. Jag sa till dem jag ville 2 pojkar och en flicka. Jag tog en gång en caben drive-in film. Filmen kostade mig $ 95.
		-- Steven Wright

%
Jag hade inga skor och jag tyckte synd själv. Sen träffade jag en man som inte hade några fötter,så jag tog hans skor.
		-- Dave Barry

%
Jag hatar när min fot somnar under dagen orsak som innebärdet kommer att vara uppe hela natten.
		-- Steven Wright

%
Jag har en låda med telefonen ringer under min säng. När jag får ensam, jagöppna upp lite, och jag får ett telefonsamtal. En dag tappade jagrutan över hela golvet. Telefonen skulle inte sluta ringa. Jag var tvungen att fådet frånkopplad. Så jag fick en ny telefon. Jag hade inte mycket pengar, så jagvar tvungen att få en oregelbunden. Det har inte en fem. Jag sprang in en vänmin på gatan häromdagen. Han sade varför inte ge mig enring upp. Jag sa att jag kan inte ringa alla jag vill längre, min telefonhar inte en fem. Han frågade hur länge det hade varit så. Jag sa att jagvisste inte - min kalender har inga sjuor.
		-- Steven Wright

%
Jag har en hund; Jag döpte honom stanna. Så när jag skulle gå att ringa honom, skulle jag säga, "Här,Stanna här ... ", men han fick klokt att det. Nu när jag ringer honom han ignorerar migoch bara håller på att skriva.
		-- Steven Wright

%
Jag har en vän vars en miljardär. Han uppfann Cliff anteckningar. NärJag frågade honom hur han fick en sådan bra idé sade han, "Jo jag först ...Jag bara ... att göra en lång historia kort ... "
		-- Steven Wright

%
Jag har en hobby. Jag har världens största samling av snäckor. jag behållerdet utspridda på stränder över hela världen. Kanske har du sett en del av det.
		-- Steven Wright

%
Jag har en karta över USA. Det är faktisk storlek. Jag tillbringade förra sommarenvika den. Folk frågar mig där jag bor, och jag säger, "E6".
		-- Steven Wright

%
Jag har ett stenparti. Förra veckan tre av dem dog.
		-- Richard Diran

%
Jag har en switch i min lägenhet som inte gör någonting. varje gångi en medan jag slår på och av. På och av. På och av. En dag jagfick ett samtal från en kvinna i Frankrike som sa "Sluta!"
		-- Steven Wright

%
Jag har en existentiell karta. Det har "Du är här" skrivet över det hela.
		-- Steven Wright

%
Jag kom precis ut från sjukhuset efter en hastighet läsning olycka.Jag träffade ett bokmärke.
		-- Steven Wright

%
Jag vet svaret! Svaret ligger i hjärtat av hela mänskligheten!Svaret är tolv? Jag tror jag är fel byggnaden.
		-- Charles Schulz

%
Jag ser på livet som kryssning chef på Titanic. Jag kan inte fådär, men jag kommer första klass.
		-- Art Buchwald

%
"Jag älskar lördag morgon tecknad film,! Detta är vad klassiska humor vadunderhållning handlar om ... Idioter, sprängämnen och fallande städ. "
		-- Calvin and Hobbes, Bill Watterson

%
Jag träffade min senaste flickvän i ett varuhus. Hon såg påkläder, och jag satte Slinkys på rulltrappor.
		-- Steven Wright

%
Jag glömmer aldrig ett ansikte, men i ditt fall ska jag göra ett undantag.
		-- Groucho Marx

%
Jag hällde fläckborttagningsmedel på min hund. Nu är han borta.
		-- Steven Wright

%
Jag satte kontaktlinser i hundens ögon. De hade lite bilder på katterpå dem. Då jag tog en ut och han sprang runt i cirklar.
		-- Steven Wright

%
Jag satte snabbkaffe i en mikrovågsugn och nästan gick tillbaka i tiden.
		-- Steven Wright

%
"Jag sa att jag hoppas att det är en bra part", säger Galder, högt."Just nu är det", säger Döden levelly. "Jag tror att det kan gåDOWNHILL mycket snabbt vid midnatt. "	"Varför?""Det var då de tror att jag ska ta min mask OFF."
		-- Terry Pratchett, "The Light Fantastic"

%
Jag såg en subliminal reklam verkställande, men bara för en sekund.
		-- Steven Wright

%
Jag borde ha varit ett land-western sångare. När allt kommer omkring, jag är äldre ände flesta västländer.
		-- George Burns

%
Jag sålde mina memoarer mitt kärleksliv till Parker Brothers - de skaatt göra ett spel av det.
		-- Woody Allen

%
Jag stannade upp hela natten spela poker med tarotkort. Jag fick en fullständighus och fyra personer dog.
		-- Steven Wright

%
Jag föreslår att du hitta din barrel utanför ditt hus, så det kommer inte att göra alltförmycket skada om det börjar brinna eller exploderar. Först bestämma vilkariktning din badtunna bör möta maximal solenergi. efter myckettrial and error, har jag funnit att den bästa riktningen för en badtunna införär uppe.
		-- Dave Barry, "The Taming of the Screw"

%
Jag säger ya, spel aldrig överens med mig. Förra veckan åkte jag till bananoch de sköt min häst med öppningen pistol.Tja, så sent som förra veckan var jag på en kinesisk restaurang och när jag öppnade minlyckokaka Jag hittade killen check sitter vid bordet bredvid. Jag sade,"Hej, kompis, jag fick din check", sade han, "Tack."
		-- Rodney Dangerfield

%
Jag tror att vi är alla bozos på denna buss.
		-- Firesign Theatre

%
Jag trodde att det var något skumt butler. Förmodligen en Fiskarna,arbetar för skala.
		-- Firesign Theatre, "The Further Adventures of Nick Danger"

%
Jag tog en kurs i läshastighet och kunde läsa Krig och fred itjugo minuter.Det handlar om Ryssland.
		-- Woody Allen

%
Jag vände luftkonditioneringsapparater tvärtom, och det blev kallt ut.Meterolog säger "Jag förstår inte det. Jag skulle vara 80grader idag, "och jag sa" Oj. "I mitt hus på taken jag har målningar av rummen ovan ... såJag har aldrig gå upp.Jag har precis köpt en mikrovågsugn spis ... Du kan tillbringa en kväll iframför den på bara åtta minuter.
		-- Steven Wright

%
Jag brukade bo i ett hus vid motorvägen. När jag gick var som helst, hade jagatt gå 65 MPH i slutet av min uppfart.Jag ersatte strålkastarna i min bil med stroboskopljus. Nu ser det utsom jag är den enda rörliga.Jag drogs över för fortkörning i dag. Officeren sade, "Vet du intehastighetsbegränsningen är 55 miles i timmen? "Och jag sa:" Ja, men jag skulle inteatt vara ute så länge. "Jag satte en ny motor i min bil, men inte ta den gamla ut. Numin bil går 500 miles i timmen.
		-- Steven Wright

%
Jag brukade arbeta i en brandpost fabrik. Du kan inte parkera någonstans näraplatsen.
		-- Steven Wright

%
Jag var på denna restaurang. Tecknet sade "Frukost som helst." Så jagbeordrade French Toast i Rennaissance.
		-- Steven Wright

%
"Jag var berusad i går kväll, kröp hem över gräsmattan. Av en slump Isätta nyckeln bil i dörrlåset. Huset startas. Så jag tänktevad fan, och körde runt kvarteret några gånger. Jag trodde jagbör gå parkera den i mitten av motorvägen och skrika åt alla attfå av min uppfart. "
		-- Steven Wright

%
Jag var i en bar och jag gick upp till en vacker kvinna och sade, "Bor durunt här ofta? "Hon sa," Du bär två olika färger strumpor. "Jag sa: "Ja, men för mig är de samma, eftersom jag går tjocklek."Hon sade, "Hur mår du?" Och jag sa: "Du vet när du sitter på enstol och du luta sig tillbaka så att du bara på två ben och du lutar alltför långt sådu nästan falla men i sista sekunden du fånga dig själv? Det känns somatt hela tiden ... "
		-- Steven Wright, "Gentlemen's Quarterly"

%
Jag var i Vegas förra veckan. Jag var vid roulettebordet, som har en långargument om vad jag ansåg ett udda tal.
		-- Steven Wright

%
Jag var det bästa jag någonsin haft.
		-- Woody Allen

%
"Jag gick in i en lanthandel, och de skulle inte sälja mig något speciellt".
		-- Steven Wright

%
"Jag gick till en anställningsintervju häromdagen frågade killen mig om jag hade någonfrågor, sa jag ja, bara ett, om du befinner dig i en bil färdas påljusets hastighet och du förvandla dina strålkastarna på, gör vad som helst hända?Han sade att han inte kunde svara på det, sa jag ledsen, men jag kunde inte arbetaför honom då.
		-- Steven Wright

%
"Jag gick till museet där de hade alla huvuden och armar frånstatyer som finns i alla andra museer. "
		-- Steven Wright

%
Jag vaknade i morse och upptäckte att allt i min lägenhethade stulits och ersatts med en exakt kopia. Jag sa till min rumskamrat,"Är inte detta fantastiskt? Allt i lägenheten har blivit stulen ochersättas med en exakt kopia. "Han sa," Jag vet att du? "
		-- Steven Wright

%
Jag arbetade i en hälsokostaffär gång. En kille kom in och frågade mig,"Om jag smälta torris, kan jag ta ett bad utan att bli blöt?"
		-- Steven Wright

%
Jag skulle hästpiska dig om jag hade en häst.
		-- Groucho Marx

%
Jag vill bli BEGRAVD indisk stil, där de sätter du upp på en hög rack,ovan jord. På så sätt kan du träffas av meteoriter och inte ensKänn det.
		-- Jack Handey, The New Mexican, 1988.

%
Jag skulle aldrig gå med i någon klubb som skulle ha sådana som mig som medlem.
		-- Groucho Marx

%
Jag kommer att vara bekväm på soffan. Kända sista ord.
		-- Lenny Bruce

%
Jag ska till Boston för att träffa min läkare. Han är en mycket sjuk människa.
		-- Fred Allen

%
Jag kommer att ge min psykoanalytiker ytterligare ett år, då kommer jag att Lourdes.
		-- Woody Allen

%
Jag kommer att leva för evigt, eller dö försöka!
		-- Spider Robinson

%
Jag är inte rädd för döden - Jag vill bara inte att vara där när det händer.
		-- Woody Allen

%
Jag har haft en helt underbar kväll. Men det var inte det.
		-- Groucho Marx

%
Om Gud hade velat att vi ska vara oroliga för den svåra situationen för de paddor, skulle hanhar gjort dem söt och lurviga.
		-- Dave Barry

%
Om bara Dionysos levde! Var skulle han äta?
		-- Woody Allen

%
Om bara Gud skulle ge mig några tydliga tecken! Som att göra en stor insättningi mitt namn på en schweizisk bank.
		-- Woody Allen, "Without Feathers"

%
Om du bor till en ålder av ett hundra du har det gjort eftersom mycket fåmänniskor dör förbi ålder av hundra.
		-- George Burns

%
Om du kastar en nyårsfest, skulle det värsta som du kan göra varaatt kasta typ av parti där dina gäster vaknar upp idag, och ringa dig för attsäger att de hade en trevlig tid. Nu kommer du att förväntas att kasta en annan partnästa år.Vad du bör göra är att kasta den typ av parti där gästen vaknaupp flera dagar från och med nu och kalla sina advokater att ta reda på om de har varitåtalade för någonting. Du vill att dina gäster att vara så angelägen att undvika enupprepning av ert parti att de omedelbart börja planera parter om derasäger, ett år i förväg, bara för att hindra dig från att ha en annan ...Om ert parti är framgångsrik, kommer polisen knackar på din dörr,såvida ert parti är mycket framgångsrik i vilket fall de kommer att LOB tårgasgenom ditt vardagsrum fönster. Som värd, är ditt jobb att se till attde inte gripa någon. Eller om de är döda uppsättning på arrestera någon,ditt jobb är att se till att det inte är du ...
		-- Dave Barry

%
Om du vill göra Gud skratta, berätta om dina planer.
		-- Woody Allen

%
Om du har gjort sex omöjliga saker före frukost, varför inte avrunda detmed middag på Milliway, restaurangen vid slutet av universum?
		-- Douglas Adams, "The Restaurant at the End of the Universe"

%
I Amerika idag ... vi har Woody Allen, vars humor har blivit såsofistikerade att ingen blir det något mer utom Mia Farrow. Alla somtror Mia Farrow ska gå tillbaka till att göra filmer där djävulen får hennegravid och Woody Allen borde gå tillbaka till att klä upp som en mänsklig spermie,du höja dina händer. Tack.
		-- Dave Barry, "Why Humor is Funny"

%
I som en dimwit, ut som ett ljus.
		-- Pogo

%
Är det konstigt här, eller är det bara jag?
		-- Steven Wright

%
Det är en viktig och populär faktum att saker och ting är inte alltid vadde verkar. Till exempel, på planeten jorden, mannen hade alltid antagitatt han var mer intelligent än delfiner eftersom han hade uppnått såmycket - hjulet, New York, krig och så vidare - medan alla delfinerhade någonsin gjort var muck om i vatten med en bra tid. Menomvänt hade delfiner alltid trott att de var långt merintelligent än människan - för exakt samma skäl.Egendomligt nog hade delfiner länge känt av den överhängandeförstörelse av planeten jorden och gjort många försök attalert mänskligheten till faran; men de flesta av deras kommunikation varmisstolkas ...
		-- Douglas Adams "The Hitchhikers' Guide To The Galaxy"

%
Det är omöjligt att uppleva en död objektivt och fortfarande bära en melodi.
		-- Woody Allen

%
Det är inte nödvändigt att ha släktingar i Kansas City för att varaolycklig.
		-- Groucho Marx

%
Det såg ut som något som liknar vit marmor, somförmodligen vad det var: något som liknar vit marmor.
		-- Douglas Adams, "The Hitchhikers Guide to the Galaxy"

%
Det är en liten värld, men jag skulle inte ha att måla den.
		-- Steven Wright

%
Det är svårt att få elfenben i Afrika, men i Alabama Tuscaloosa.
		-- Groucho Marx

%
Det är inte att jag är rädd för att dö. Jag vill bara inte att vara där när det händer.
		-- Woody Allen

%
I går kväll strömmen gick ut. Bra min kamera hade en blixt ....Grannarna trodde att det var blixten i mitt hus, så de kallade polisen.
		-- Steven Wright

%
Förra året körde vi över hela landet ... Vi bytte på driv ...varje halv mil. Vi hade ett kassettband att lyssna på hela resan.Jag minns inte vad det var.
		-- Steven Wright

%
Livet är uppdelad i den fruktansvärda och olycklig.
		-- Woody Allen, "Annie Hall"

%
Livet går till spillo på de levande.
		-- The Restaurant at the End of the Universe.

%
Precis som ni, jag ofta hemsökt av djupgående frågor som rör människansplats i systemet av saker. Här är några:Q - Finns det liv efter döden?A - Definitivt. Jag talar av egen erfarenhet här. på NewNyårsafton, 1970, drack jag en hel kanna av en drink som heter "Black Russian",sedan kröp ut på gräsmattan och dog inom några minuter, vilket varbra med mig eftersom jag hade insett att om jag hade levt jag skulle habringade resten av mitt liv i klorna på de otroligt smärtsamthuvudvärk. Tack vare miraklet med modern apelsinjuice, jag kom tillbakatill livet flera dagar senare, men under tiden jag var definitivt död. jagantar att min huvudsakliga intryck av livet efter detta är att det är inte så illa så längesom du håller TV tackade och inte försöka äta någon fast föda.
		-- Dave Barry

%
Man 1: Fråga mig vad det viktigaste om att berätta en bra skämt är.Man 2: OK, vad är det mest impo -Man 1: ______ timing!
		-- Dave Barry

%
"Många har sett Topaxci, Gud Röda svamp, och de tjänarnamn på shaman, "säger han. Några har sett Skelde, andan i rök, ochDe kallas trollkarlar. Några har haft förmånen att se Umcherrel, densjäl i skogen, och de är kända som ande mästare. Men ingen harsett en låda med hundratals ben som såg på dem utan ögon, och deär kända som idio-- "Avbrottet orsakades av en plötslig skrikande ljud och en uppsjösnö och gnistor som blåste elden över mörka hut; det fanns en kortdimsyn och sedan den motsatta väggen sprängdes undan ochuppenbarelse försvunnit.Det blev en lång tystnad. Sedan en något kortare tystnad. Sedanden gamla shamanen sade noggrant, "Du har inte bara se två män gå igenomupp och ner på en kvast, skrika och skriker på varandra, eller hur? "Pojken såg på honom levelly. "Absolut inte", sade han.Den gamle mannen drog en suck av lättnad. "Tack och lov för det," hansa. "Inte heller jag."
		-- Terry Pratchett, "The Light Fantastic"

%
Många år sedan under en period som vanligtvis känner som nästa fredag ​​eftermiddag,bodde en kung som var mycket dyster på tisdag morgon eftersom hanvar så Sad tänkande om hur olycklig han hade varit på måndag och hurhelt Sorglig han skulle vara på onsdag ....
		-- Walt Kelly

%
Min bror skickade mig ett vykort häromdagen med denna stora satellitbildav hela jorden på den. På baksidan det sade: "Önskar du var här".
		-- Steven Wright

%
Min vän har en baby. Jag skriver ner alla ljud han gör såsenare jag kan fråga honom vad han menade.
		-- Steven Wright

%
Mina vänner, jag är här för att berätta om den wonderous kontinenten kallasAfrika. Väl vi lämnade New York berusad och tidigt på morgonen den 31 februari.Vi var 15 dagar på vattnet, och tre på båten när vi äntligen kom iAfrika. Vid vår ankomst vi omedelbart inrätta ett rigoröst schema: Upp till06:00, frukost, och tillbaka i sängen med 07:00. Ganska snart var vi tillbaka i sängen med06:30. Nu Afrika är full av stora spelet. Den första dagen jag sköt två dollar. Den därvar det största spelet som vi hade. Afrika är primerally bebos av Elks, Mooseoch riddarna av Pithiests.Älgarna lever upp i bergen och komma ner en gång om året för sinårliga konventioner. Och du bör se dem samlades runt vattenhålet,som de lämnar omedelbart när de upptäcker att det är full av vatten. Devar inte ute efter ett vattenhål. De letade efter en alck hål.En morgon jag sköt en elefant i min pyjamas, hur han fick i minpyjamas, jag vet inte. Sedan försökte vi att ta bort betar. Det är en tufford att säga, betar. Som sagt vi försökte ta bort beta, men de varinbäddad så hårt vi inte kunde få ut dem. Men i Alabama Tuscaloosa,men det är helt Irrelephant vad jag sade.Vi tog några bilder av de infödda flickor, men de var inte utvecklats.Så vi kommer tillbaka om några år ...
		-- Julius H. Marx [Groucho]

%
Nietzsche säger att vi kommer att leva samma liv, om och om igen.Gud - Jag måste sitta igenom isen Capades igen.
		-- Woody Allen, "Hannah and Her Sisters"

%
Nirvana? Det är den plats där de krafter som och deras vänner umgås.
		-- Zonker Harris

%
Ingen förväntar sig den spanska inkvisitionen!
		-- Zonker Harris

%
Nu är det dags för alla goda män att komma till.
		-- Walt Kelly

%
Uppenbarligen föremål för döden var i luften, men mer som någotundvikas än harped på.Möjligen den fasa som Zaphod upplevde vid tanken på att varaåterförenas med sina avlidna släktingar ledde till tanken att de kanbara känner på samma sätt om honom och, vad mer, kunna göra någotom att hjälpa att skjuta denna återförening.
		-- Douglas Adams

%
Man behöver inte ha ett sinne för humor. Det har du.
		-- Larry Gelbart

%
Utanför en hund, är en bok människans bästa vän. Inne i en hund är det ocksåmörk att läsa.
		-- Groucho Marx

%
Vitsar är lite "spelar på orden" att en viss typ av person som älskar attvåren på dig och sedan titta på dig i en viss självbelåten sätt atttyder på att han tror att du måste tro att han är den i särklass smartasteperson på jorden nu att Benjamin Franklin är död, när i själva verket vad dutänker är att om denna person någonsin hamnar i en livbåt, den andrapassagerarna kasta honom överbord i slutet av den första dagen, även om dehar gott om mat och vatten.
		-- Dave Barry, "Why Humor is Funny"

%
"Just nu jag har minnesförlust och deja vu samtidigt."
		-- Steven Wright

%
Rincewind bildade en mental bild av någon underlig enhet som bor i ett slottgjord av tänder. Det var typ av mental bild du försökte glömma.Utan framgång.
		-- Terry Pratchett, "The Light Fantastic"

%
Romeo inte bilked i en dag.
		-- Walt Kelly, "Ten Ever-Lovin' Blue-Eyed Years With Pogo"

%
Hajar är lika tuff som de fotbollsfans som tar sina skjortor avunder spel i Chicago i januari bara mer intelligent.Tonåring bör veta "
		-- Dave Barry, "Sex and the Single Amoeba: What Every

%
Dyka upp är 80% av livet.
		-- Woody Allen

%
Några av er ... kanske har beslutat att i år, kommer du att firaden gammaldags sätt, med din familj sitter runt strängtranbär och utbyta ödmjuka, handgjorda presenter, som på "The Waltons".Tja, kan du glömma det. Om alla drog den typen av subversiva stunt,ekonomin skulle kollapsa under natten. Regeringen skulle behövaingripa: det skulle bilda ett kabinett-nivå Institutionen för Holiday julklapparna,vilket skulle spendera miljarder och åter miljarder av skattepengar för att köpa Barbiedockoroch elektroniska spel, som det skulle falla på befolkningen från flygvapnetjets, döda och lemlästa tusentals. Så, till gagn för nationen, dubör gå tillsammans med Holiday Program. Detta innebär att du ska få en storsumma pengar och gå till ett köpcentrum.
		-- Dave Barry, "Christmas Shopping: A Survivor's Guide"

%
Ibland skönheten i världen är så överväldigande, jag vill bara att kastatillbaka mitt huvud och gurgla. Bara gurgla och gurgla och jag bryr mig inte som hörmig eftersom jag är vacker.
		-- Jack Handey, The New Mexican, 1988.

%
Tack och lov modern bekvämlighet är ett minne avlägsen framtid.
		-- Pogo, by Walt Kelly

%
Den grundläggande idén bakom varuhus är att de är mer praktiskt än städer.Städer innehåller gator, som är farliga och trångt och svårt attpark i. varuhus, å andra sidan, har parkeringsplatser, som också ärfarlig och trångt och svårt att parkera på, men - här är den storaskillnad - i köpcentret parkeringsplatser, det finns inga regler. Du är tillåtet attgör något. Du kan köra så fort du vill ha i någon riktning du vill.Jag var en gång kör i ett köpcentrum parkeringsplats när min bil träffades av en pickuplastbil drivs bakåt av en knäböj man med en tatuering som sa "Charlie"på hans underarm, som kom ut och förklarade för mig, i detalj, varförolyckan var mitt fel, hans resonemang är att han var våldsam och muskulös,medan jag var varken. Denna typ av resonemang är juridiskt giltigt i köpcentretparkeringsplatser.
		-- Dave Barry, "Christmas Shopping: A Survivor's Guide"

%
Det bästa botemedlet mot sömnlöshet är att få mycket sömn.
		-- W. C. Fields

%
Det bästa sättet att göra upp eld med två pinnar är att se till att en av demär en match.
		-- Will Rogers

%
Buffalo är inte lika farligt som alla gör honom att vara.Statistiken visar att fler amerikaner i USA dödas ibilolyckor än dödas av buffel.
		-- Art Buchwald

%
Den stora språng i valen upp nedgången av Niagara är uppskattade, av allasom har sett den, som en av de finaste glasögon i naturen.
		-- Benjamin Franklin.

%
Liftarens guide till galaxen har några saker att säga omföremål för handdukar.Viktigast har en handduk enorm psykologisk värde. Förnågon anledning, om en icke-liftare upptäcker att en liftare har sin handdukmed honom, kommer han automatiskt anta att han är också i besittning av entandborste, tvättlapp, kolv, gnat spray, rymddräkt, etc., etc. Dessutom,den icke-liftare kommer sedan glatt låna ut liftare någon av dessa ellerett dussin andra objekt som han kan ha "förlorat". När allt kommer omkring, som någon människa kanhitch längden och bredden av Galaxy, kämpa mot fruktansvärda odds,vinna igenom och fortfarande vet var hans handduk är, är uppenbarligen en man att vararäkna med.
		-- Douglas Adams, "The Hitchhiker's Guide to the Galaxy"

%
Den andra dagen jag ... eh, nej, det var inte jag.
		-- Steven Wright

%
"Pyramiden öppnar!"	"Vilken?""Den med allt större hål i det!"När när du inte någonstans alls "
		-- Firesign Theater, "How Can You Be In Two Places At

%
De tre stora typ av verktyg* Verktyg för hittings saker att göra dem lös eller att skärpa dem ellerjar sina många komplexa, sofistikerade elektriska delar på ett sådantsätt att de fungerar perfekt. (Detta är dina hammare, spikklubbor,klubbor och batonger.)* Verktyg som, om den tappas på rätt sätt, kan tränga foten. (Sylar)* Verktyg som ingen någonsin skulle använda eftersom den potentiella faran är långtstörre än värdet av ett projekt som eventuellt skulle kunna leda till.(Motorsågar, borrmaskiner, kraft häftapparater, någon form av verktyg som användernågon form av makt mer avancerad än ficklampa batterier.)
		-- Dave Barry, "The Taming of the Screw"

%
Det kommer en tid i angelägenheter en man när han måste ta tjureni svansen och möta situationen.
		-- W. C. Fields

%
Det finns inget enkelt snabbt sätt ut, vi ska ha för att leva genom vårhela livet, vinna, förlora eller rita.
		-- Walt Kelly

%
Det finns så mycket plast i denna kultur som vinyl leopardskinn ärbli en hotad syntetiska.
		-- Lily Tomlin

%
Det kommer att bli bättre trots våra ansträngningar för att förbättra dem.
		-- Will Rogers

%
Detta land är fullt av byxor!detta land är fullt av mausergevär!Och Pussycats att äta dem när solen går ner!
		-- Firesign Theater

%
Tid är en illusion, lunchtid dubbelt så.
		-- The Hitchhiker's Guide to the Galaxy

%
Synd att du inte kan köpa en voodoo världen så att du kan göra jorden snurrariktigt snabbt och missfoster ut alla.
		-- Jack Handey, The New Mexican, 1988.

%
Tjugo procent av Zero är bättre än ingenting.
		-- Walt Kelly

%
Vi har mött fienden, och han är oss.
		-- Walt Kelly

%
Vi konfronteras med oöverstigliga möjligheter.
		-- Walt Kelly, "Pogo"

%
Vad händer om allt är en illusion och ingenting existerar? I så fall, jagdefinitivt betalat för mycket för min matta.
		-- Woody Allen, "Without Feathers"

%
Vad händer om ingenting existerar och vi är alla i någons dröm? Eller vad värre är,vad händer om bara att fett killen i den tredje raden finns?
		-- Woody Allen, "Without Feathers"

%
Vad är komedi? Komedi är konsten att få människor att skratta utan att göradem spy.
		-- Steve Martin

%
	"Vad ska vi göra?" sade Twoflower."Panic?" sade Rincewind förhoppningsvis. Han höll alltid att panik vardet bästa sättet att överleva; tillbaka i gamla tider, hans teori gick, människorinför hungriga sabretoothed tigrar kunde delas mycket enkelt inde som panik och de som stod där säger "Vad en magnifikkräk! "och" Här fitta. "
		-- Terry Pratchett, "The Light Fantastic"

%
Vad är ett annat ord för "synonymordbok"?
		-- Steven Wright

%
När jag var över gränsen till Kanada, frågade de omJag hade några skjutvapen med mig. Jag sa: "Ja, vad behöver du?"
		-- Steven Wright

%
När jag var liten, gick jag in i en djuraffär och de frågade hur stor jag skulle få.
		-- Rodney Dangerfield

%
När jag vaknade i morse, frågade min flickvän om jag hade sovit gott.Jag sa: "Nej, jag gjorde några misstag."
		-- Steven Wright

%
Där humor är oroad finns det inga normer - ingen kan säga vadär bra eller dåligt, men du kan vara säker på att alla kommer.
		-- John Kenneth Galbraith

%
Varför är alfabetet i den ordningen? Är det på grund av den låten?
		-- Steven Wright

%
Will Rogers aldrig träffat dig.
		-- Steven Wright

%
Winny och jag bodde i ett hus som körde på statisk elektricitet ...Om du vill köra mixer, var du tvungen att gnugga ballonger påhuvud ... om du vill laga mat, var du tvungen att dra bort en tröja riktigt snabbt ...
		-- Steven Wright

%
Vill du * ______ verkligen * vill komma på en non-stop flyg?
		-- George Carlin

%
Du kan inte få allt. Var skulle du säga?
		-- Steven Wright

%
"Du vet, det är ibland så här när jag fångade i en Vogonluftsluss med en man från Betelgeuse och på väg att dö av kvävning irymden som jag önskar verkligen att jag hade lyssnat på vad min mamma berättadenär jag var ung!""Varför, vad hon sa?""Jag vet inte, jag lyssnade inte."
		-- Douglas Adams, "The Hitchhiker's Guide to the Galaxy"

%
Du kanske redan vara en förlorare.
		-- Form letter received by Rodney Dangerfield.

%
Du skulle bättre slå det. Du kan lämna i en taxi. Om du inte kan få en taxi, dukan lämna in en huff. Om det är för tidigt, kan du lämna in en minut och en huff.
		-- Groucho Marx

%
Du är ett bra exempel på varför vissa djur äter sina ungar.Ja, just det. Jag minns min första öl.När din IQ stiger till 28, sälja.
		-- Professor Irwin Corey to a heckler

%
FORTUNE Random citerar match spel 75, NO. 1: Gene Rayburn: Vi skulle vilja avsluta med en tanke för dagen, vänner ---               något ...      Någon: (avbryter) Uh-oh Gene Rayburn: ... kärnfulla, full av visdom --- och vi uppmanar Poet               Laureate, Nipsey RussellNipsey Russell: Ungdomarna är mycket annorlunda i dag, och det finns               ett säkert sätt att veta: Barn används för att fråga var de kom               från, nu kommer de att tala om var du kan gå.          Alla: (skratt)
		-- Professor Irwin Corey to a heckler

%
