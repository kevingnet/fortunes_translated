17 Rule of Friendship:En vän kommer att avstå från att berätta att han plockade upp samma mängdliv försäkringsskydd du gjorde för halva priset när din ärej annullerbara.
		-- Esquire, May 1977

%
186,282 miles per sekund:Det är inte bara en bra idé, det är lagen!
		-- Esquire, May 1977

%
18 Rule of Friendship:        En vän låter dig hålla stegen medan han går upp på taket        att installera din nya antenn, som är den största son-of-a-tik du        någonsin sett.
		-- Esquire, May 1977

%
2180, US History fråga:Vad 20th Century USA: s president var nästan inför riksrätt och vadkontor gjorde han senare hålla?
		-- Esquire, May 1977

%
3rd lag Computing:Allt som kan gå wrförmögenhet: Segmente överträdelse - Kärna dumpas
		-- Esquire, May 1977

%
667:Grannen av odjuret.
		-- Esquire, May 1977

%
Ett hypotetiskt paradox:Vad skulle hända i en strid mellan en Enterprise säkerhetsgruppsom alltid dödas strax efter visas och en trupp av ImperialStormtroopers, som inte kan slå den breda sidan av en planet?
		-- Tom Galloway

%
En lag Datorprogrammering:Gör det möjligt för programmerare att skriva på engelskaoch du kommer att tycka att programmerare inte kan skriva på engelska.
		-- Tom Galloway

%
En musiker, konstnär, arkitekt:den man eller kvinna som inte är en av dessa är inte en kristen.
		-- William Blake

%
En ny koan:Om du har några glass, kommer jag ge det till dig.Om du inte har någon glass, kommer jag att ta det ifrån dig.Det är en glass koan.
		-- William Blake

%
Abbotts råden:(1) Om du måste fråga, du är inte rätt att få veta.(2) Om du inte gillar svaret, du skulle inte ha ställt frågan.
		-- Charles Abbot, dean, University of Virginia

%
Frånvarande, adj .:Utsätts för angrepp av vänner och bekanta; förtalas; förtalad.
		-- Charles Abbot, dean, University of Virginia

%
Frånvarande, n .:En person med en inkomst som har haft eftertanke för att ta bortsig från området för exactionen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Abstainer, n .:En svag person som ger efter för frestelsen att förneka sig själv ennöje.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Absurditet, n .:Ett uttalande eller övertygelse uppenbart oförenligt med en egen uppfattning.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Akademi:En modern skola där fotboll lärs ut.Inleda:En ålderdomlig skola där fotboll inte lärs ut.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Acceptanstest:Ett misslyckat försök att hitta fel.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Olycka, n .:Ett tillstånd där sinnesnärvaro är bra, men avsaknaden avkroppen är bättre.
		-- Foolish Dictionary

%
Dragspel, n .:En säckpipe med veck.
		-- Foolish Dictionary

%
Noggrannhet, n .:Vice av att vara rätt
		-- Foolish Dictionary

%
Bekant, n:En person som vi känner väl tillräckligt för att låna från, men inte branog att låna ut till. En viss grad av vänskap som kallas lätt närobjektet är dålig eller oklar, och intim när han är rik eller berömd.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
ADA:Något du behöver bara veta namnet på att vara en expert iComputing. Användbar i meningar som: "Vi hade bättre utvecklaen ADA medvetande.
		-- "Datamation", January 15, 1984

%
Adler distinktion:Språket är allt som skiljer oss från de lägre djuren,och från byråkraterna.
		-- "Datamation", January 15, 1984

%
Beundran, n .:Vår artig erkännande av varandras likheter med oss.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Adore, v .:Att vörda förväntans.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Vuxen, n .:En gammal nog att veta bättre.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Reklam Regel:Skriftligen en patentmedicin annonsering, först övertygaläsare som han har sjukdomen han läser om, för det andra,att det kan botas.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Eftermiddag, n .:Den del av dagen vi spenderar oroa dig för hur vi slösat bort på morgonen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ålder, n .:Denna period i livet där vi förening för laster som vifortfarande vårda genom smäda dem som vi inte längre har företaget	att begå.
		-- Ambrose Bierce

%
Agnes lag:Nästan allt i livet är lättare att komma in än ut ur.
		-- Ambrose Bierce

%
Air Force Inertia Axiom:Konsekvens är alltid lättare att försvara än korrekthet.
		-- Ambrose Bierce

%
luft, n .:En näringsrik substans som tillhandahålls av en riklig försyn förgödning av de fattiga.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Alaska:Ett förspel till "Nej"
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Albrecht lag:Sociala innovationer tenderar att nivån på minimi acceptabel välbefinnande.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Alden s lagar:(1) Ge bort babykläder och möbler är den största orsakenav graviditeten.(2) alltid vara bakgrundsbelyst.(3) Sitt ner när det är möjligt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
algoritm, n .:Trendig dans för höft programmerare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
underhållsbidrag, n:Med en ex du kan satsa på.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Allt nytt:Delar inte utbytbara med tidigare modell.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Allens Axiom:När allt annat misslyckas, läs instruktionerna.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Alliance, n .:I den internationella politiken, en förening av två tjuvar som harderas händer så djupt in i varandras ficka att de inte kanseparat plundra tredjedel.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ensam, adj .:I dåligt sällskap.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ambidextrous, adj .:Kunna plocka med samma skicklighet en högerficka eller vänster.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Tvetydighet:Talar sanning när du inte meningen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ambition, n:En overmastering önskan att bli förtalad av fiender medanlevande och gjort löjligt av vänner när död.
		-- Ambrose Bierce

%
Amoebit:Amöba / kanin kors; det kan multiplicera och dividera samtidigt.
		-- Ambrose Bierce

%
Andreas förmaning:skänka aldrig svordomar på en förare som har kränkt dig.Om du tror att hans fönster är stängda och han kan inte höra dig,det är inte och han kan.
		-- Ambrose Bierce

%
Androphobia:Rädsla för män.
		-- Ambrose Bierce

%
Smörja, v .:Att smörja en kung eller andra stora funktionär redan tillräckligthala.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Anthony lag om Force:Tvinga inte; få en större hammare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Anthony lag av Workshop:Alla verktyg när de släpps, kommer att rulla in i minst åtkomlighörnet av verkstaden.Naturlig följd:På vägen till hörnet, kommer någon tappat verktyg först slåtårna.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Antonym, n .:Motsatsen till ordet du försöker att tänka på.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Afasi:Förlust av tal i samhällsvetare när badpå fester, "Men vilken nytta är din forskning?"
		-- Ambrose Bierce, "The Devil's Dictionary"

%
aforism, n .:En kortfattad, smart uttalande.afterism, n .:En kortfattad, smart uttalande du inte tänker på förrän alltför sent.
		-- James Alexander Thom

%
Bilaga:En del av en bok, för vilken ingen ännu har upptäckt någon användning.
		-- James Alexander Thom

%
Applåder, n:Ekot av en plattityd från mynningen av en dåre.
		-- Ambrose Bierce

%
aquadextrous, adj .:Besitter förmågan att vända badkaret kran på och utanförmed tårna.
		-- Rich Hall, "Sniglets"

%
Godtyckliga system pl.n .:System om vilken inget allmänt kan sägas, spara "ingentingallmänhet kan sägas. "
		-- Rich Hall, "Sniglets"

%
Aritmetisk:En obskyr art inte längre praktiseras i världens industriländer.
		-- Rich Hall, "Sniglets"

%
bältdjur:Att ge vapen till en spansk knipa.
		-- Rich Hall, "Sniglets"

%
Rustning Axiom:Dygd är misslyckandet med att uppnå vice.
		-- Rich Hall, "Sniglets"

%
Armstrong samling lag:Om kontrollen är verkligen i posten,Det är säkerligen gjord till någon annan.
		-- Rich Hall, "Sniglets"

%
Arnolds Addendum:Allt som inte passar in i dessa kategorier orsakar cancer hos råttor.
		-- Rich Hall, "Sniglets"

%
Arnolds lagar Documentation:(1) Om det skulle existera, det gör det inte.(2) Om det existerar, är den inaktuell.(3) Endast dokumentation för onödiga program överskridertvå första lagar.
		-- Rich Hall, "Sniglets"

%
Arthur lagar Kärlek:(1) Människor som du lockas alltid tror att dupåminna dem om någon annan.(2) Den kärleksbrev du äntligen modet att skicka blirförsenade i post tillräckligt länge för att göra narr avsjälv personligen.
		-- Rich Hall, "Sniglets"

%
ASCII:Styrkoden för alla börjar programmerare och de som skullebli datorvana. Etymologiskt har termen kommit ned somen sammandragning av ofta upprepade frasen "ascii och du skall	ta emot."
		-- Robb Russon

%
Atlanta:En hel stad omgiven av en flygplats.
		-- Robb Russon

%
Auktion:En gyp bort den gamla block.
		-- Robb Russon

%
audiophile, n:Någon som lyssnar till utrustningen i stället för musiken.
		-- Robb Russon

%
Äkta:Otvivelaktigt sant, i någon mening.
		-- Robb Russon

%
Automobile, n .:En fyrhjuligt fordon som går upp kullar och ned fotgängare.
		-- Robb Russon

%
Ungkarl:En kille som är rotlösa och fästmö fritt.
		-- Robb Russon

%
Ungkarl:En man som jagar kvinnor och aldrig Mrs en.
		-- Robb Russon

%
Bakåt konditionering:Att sätta saliv i en hunds mun i ett försök att göra en klocka ring.
		-- Robb Russon

%
Bagbiter:1. n .; Utrustning eller program som misslyckas, oftast intermittent. 2.adj .: misslyckas hårdvara eller mjukvara. "Detta bagbiting systemet inte kommer att låta mig fåav Spacewar "Användning: vägrenar på obscenitet Grammatically avskiljas, en..kan tala om "bita påsen". Synonymer: förlorare, förlora, KRETINISK,BLETCHEROUS, BARFUCIOUS, Chomper, chomping.
		-- Robb Russon

%
Bagdikian Observations:Försöker vara en första klassens reporter på den genomsnittliga amerikanska tidningenär som att försöka spela Bachs "Matteuspassionen" på en ukelele.
		-- Robb Russon

%
Baker första lag av Federal geometri:Ett block bidrag är en fast massa pengar omgiven på alla sidor avguvernörer.
		-- Robb Russon

%
Ballistophobia:Rädsla för kulor;Otophobia:Rädsla för att öppna sina ögon.Peccatophobia:Rädsla för att synda.Taphephobia:Rädsla för att bli levande begravda.Sitophobia:Rädsla för livsmedel.Trichophobbia:Rädsla för hår.Vestiphobia:Rädsla för kläder.
		-- Robb Russon

%
Banacek artonde polska ordspråket:Flodhästen har ingen sting, men den vise mannen skulle snarare vara satt påav bi.
		-- Robb Russon

%
Banectomy, n .:Avlägsnandet av blåmärken på en banan.
		-- Rich Hall, "Sniglets"

%
Barach härskar:En alkoholist är en person som dricker mer än sin egen läkare.
		-- Rich Hall, "Sniglets"

%
Barbara arbetsordning bitter erfarenhet:(1) När du tömmer en låda för sina kläderoch en hylla för sina toalettartiklar, avslutar relationen.(2) När du äntligen köpa ganska stillaatt fortsätta korrespondens, stannar han skriva.
		-- Rich Hall, "Sniglets"

%
Barkers Bevis:Korrekturläsning är effektivare efter offentliggörandet.
		-- Rich Hall, "Sniglets"

%
Barometer, n .:En sinnrik instrument som visar vilken typ av väder vi	har.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Barth distinktion:Det finns två typer av människor: de som delar in människor i tvåtyper, och de som inte gör det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Baruchs Observation:Om allt du har är en hammare, allt ser ut som en spik.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Grundläggande definitioner of Science:Om det är grönt eller wiggles, det är biologi.Om det stinker, det är kemi.Om det inte fungerar, är det fysik.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
BASIC, n .:Ett programmeringsspråk. Relaterade till vissa sociala sjukdomar iatt de som har det kommer inte att erkänna det i artigt företag.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bathquake, n .:Den våldsamma skalv som skramlar hela huset när vattnetkran är påslagen till en viss punkt.
		-- Rich Hall, "Sniglets"

%
Strid, n .:En metod för obundet med tänderna en politisk knut somkommer inte att ge på tungan.
		-- Ambrose Bierce

%
Skönhet, n .:Kraften med vilken en kvinna charm en vän och skrämmer en make.
		-- Ambrose Bierce

%
Skönhet:Vad som finns i ögat när du har ett bi i handen.
		-- Ambrose Bierce

%
Begathon, n .:En flera dagar evenemang på den statliga televisionen, som används för att samla in pengar sådu kommer inte att titta på reklam.
		-- Ambrose Bierce

%
Beifeld princip:Sannolikheten för en ung man möte en önskvärd och mottagligunga kvinnliga ökar med pyramid progression när hanär redan i sällskap med (1) ett datum, (2) hans fru, (3) ensnyggare och rikare manliga vän.
		-- R. Beifeld

%
tro, n:Något du inte tror.
		-- R. Beifeld

%
Bennetts lagar trädgårdsnäring:(1) Husen är för människor att leva i.(2) Gardens är för växter att leva i.(3) Det finns inget sådant som en krukväxt.
		-- R. Beifeld

%
Benson Dogma:ASCII är vår gud, och Unix är hans vinst.
		-- R. Beifeld

%
Bershere Formel för misslyckande:Det finns bara två typer av människor som misslyckas: de somlyssna på ingen ... och de som lyssnar på alla.
		-- R. Beifeld

%
beta test, v:Att frivilligt anförtro sina uppgifter, en försörjning och sinförnuft till maskin- eller programvara avsedd för att förstöra alla tre.I tidigare dagar, var oskulder ofta väljs för betatestning vulkaner.
		-- R. Beifeld

%
Bierman lagar Kontrakt:(1) I varje dokument, kan du inte täcka alla "tänk om är".(2) Advokater stanna kvar i verksamheten att lösa alla olösta "tänk om är".(3) Varje löst "tänk om" skapar två olösta "tänk om är".
		-- R. Beifeld

%
Bilbos första lag:Du kan inte räkna vänner som alla är förpackade i fat.
		-- R. Beifeld

%
Binär, adj .:Ha förmåga att ha vänner av båda könen.
		-- R. Beifeld

%
Bing Regel:Försök inte att hejda - flytta stranden.
		-- R. Beifeld

%
Bipolär, adj .:Avser någon som har hem i Nome, Alaska, och Buffalo, New York.
		-- R. Beifeld

%
födelse, n:Den första och direst av alla katastrofer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
bit, n:En måttenhet tillämpas på färg. Tjugofyra-bitars färghänvisar till dyra $ 3 färg i motsats till den billigare 25cent, eller två-bitars, färg som använder för att vara tillgängliga för några år sedan.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bizoos, n .:De miljontals små enskilda gupp som utgör en basketboll.
		-- Rich Hall, "Sniglets"

%
blithwapping:Med hjälp av något annat än en hammare för att hamra en spik i denvägg, såsom skor, lampfötter, dörrs, etc.
		-- "Sniglets", Rich Hall & Friends

%
Bloom sjunde lag Litigation:Domarens skämt är alltid roligt.
		-- "Sniglets", Rich Hall & Friends

%
Blore rakkniv:Med tanke på ett val mellan två teorier, ta den som är roligare.
		-- "Sniglets", Rich Hall & Friends

%
Blutarsky s Axiom:Ingenting är omöjligt för den som inte kommer att ta reson.
		-- "Sniglets", Rich Hall & Friends

%
Boling postulatet:Om du känner dig bra, oroa dig inte. Du kommer över det.
		-- "Sniglets", Rich Hall & Friends

%
Bolub fjärde lag Computerdom:Projektgrupper avskyr veckolägesrapportering eftersom det sålivligt visar deras brist på framsteg.
		-- "Sniglets", Rich Hall & Friends

%
Bombeck s Rule of Medicine:Aldrig gå till en läkare vars kontor växter har dött.
		-- "Sniglets", Rich Hall & Friends

%
Boob lag:Du hittar alltid något på det sista stället du ser ut.
		-- "Sniglets", Rich Hall & Friends

%
Booker lag:Ett uns av ansökan är värt massor av abstraktion.
		-- "Sniglets", Rich Hall & Friends

%
Bore, n .:En kille som sveper upp en två minuters idé i en två-timmars ordförråd.
		-- Walter Winchell

%
Bore, n .:En person som talar när du önskar honom att lyssna.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Boren s lagar:(1) När ansvaret, fundera.(2) När du är i trubbel, delegera.(3) Om du är osäker, mumla.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
chef, n:Enligt Oxford English Dictionary, i medeltidenOrden "boss" och "fuskverk" var i stort sett synonymt med undantag av att chefen,förutom betyder "en handledare för arbetare" också inneburit "enprydnads stud. "
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bouchers Observation:Han som blåser sin egen horn alltid spelar musikflera oktaver högre än vad som ursprungligen skriven.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bower lag:Talang går där det händer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bowies Sats:Om ett experiment fungerar måste du använda fel utrustning.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
pojke, n:En brus med smuts på den.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bradleys Bromid:Om datorer blir för stark, kan vi organiseradem i en kommitté - som kommer att göra dem.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Brady första lag problemlösning:När de konfronteras med ett svårt problem, kan du lösa det merlätt genom att reducera den till frågan, "Hur skulle Lone Rangerhar hanterat detta? "
		-- Ambrose Bierce, "The Devil's Dictionary"

%
hjärna, n:Apparaten som vi tror att vi tror.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
hjärna, v: [som i "till hjärnan"]Att tillrätta rakt på sak, men inte tillspetsat; att skingra en källaav fel i en motståndare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
hjärnskadade, generalisering av "Honeywell Brain Damage" (HBD), enteoretisk sjukdom uppfanns för att förklara vissa fullkomlig cretinisms iMultics, adj:Uppenbarligen fel; KRETINISK; tokig. Det finns en implicitatt den person som ansvarar måste ha lidit hjärnskador,eftersom han / hon borde ha vetat bättre. Calling någothjärnskadade är dålig; det innebär också att det är oanvändbart.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bride, n .:En kvinna med en fin utsikt av lycka bakom henne.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
portfölj, n:En studie där juryn får tillsammans och bildar en lynchning part.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
vidsynthet, n:Resultatet av platt hög sinne ut.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Brogan s Konstant:Människor tenderar att samlas på baksidan av kyrkan ochframför bussen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
brokee, n:Någon som köper aktier på inrådan av en mäklare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Brontosaurus Princip:Organisationer kan växa snabbare än deras hjärnor kan hantera demi förhållande till sin omgivning och sin egen fysiologi: närdetta sker, de är en utrotningshotad art.
		-- Thomas K. Connellan

%
Bäck lag:Lägga arbetskraft till en sen programvaruprojekt gör det senare.
		-- Thomas K. Connellan

%
Brookes lag:Närhelst ett system blir fullständigt definierad, vissa idiotupptäcker något som antingen avskaffar systemet ellerexpanderar den till oigenkännlighet.
		-- Thomas K. Connellan

%
Bubbla minne, n .:En nedsättande term, vanligen med hänvisning till en persons intelligens.Se även "vakuumrör".
		-- Thomas K. Connellan

%
Bucy lag:Ingenting är någonsin åstadkommas genom en förnuftig människa.
		-- Thomas K. Connellan

%
Bug, n .:En aspekt av ett datorprogram som finns på grund av attprogrammerare tänkte Jumbo Jacks or optioner när han / honskrev programmet.Lyckligtvis har näst sista bugg bara rättats.
		-- Ray Simard

%
bug, n:En son till en glitch.
		-- Ray Simard

%
bug, n:En gäckande varelse som lever i ett program som gör det fel.Aktiviteten hos "felsökning", eller ta bort fel från ett program slutarnär folk tröttnar på att göra det, inte när buggar tas bort.
		-- "Datamation", January 15, 1984

%
Buggar, pl. n .:Små levande saker som små levande pojkar kasta på små levande flickor.
		-- "Datamation", January 15, 1984

%
Bildekal:Alla de delar som faller utanför denna bil är av allra finasteBritish tillverkning.
		-- "Datamation", January 15, 1984

%
Bunker förmaning:Du kan inte köpa öl; du kan bara hyra den.
		-- "Datamation", January 15, 1984

%
Burbulation:Den tvångshandling att öppna och stänga en kylskåpsdörr iett försök att fånga den innan den automatiska ljuset tänds.
		-- "Sniglets", Rich Hall & Friends

%
Bureau uppsägning, lag:När en regering byrå är planerad att fasas ut,Antalet anställda i den byrå kommer att fördubblas inom12 månader efter det att beslut fattas.
		-- "Sniglets", Rich Hall & Friends

%
byråkrati, n:En metod för att omvandla energi till fast avfall.
		-- "Sniglets", Rich Hall & Friends

%
Byråkrat, n .:En person som minskar byråkratin i sidled.
		-- J. McCabe

%
byråkrat, n:En politiker som har besittningsrätt.
		-- J. McCabe

%
Burke postulat:Allt är möjligt om du inte vet vad du talar om.Skapa inte ett problem som du har inte svaret.
		-- J. McCabe

%
Bränn Hog ​​vägningsmetod:(1) Få en perfekt symmetrisk planka och balansera det över en sågbock.(2) Placera hog på en ände på plankan.(3) Pile stenar på den andra änden tills plankan är åter perfektbalanserad.(4) antar vikten hos stenarna försiktigt.
		-- Robert Burns

%
modeord, n:Smolket i glädjebägaren av datakunskap.
		-- Robert Burns

%
byob, volym:Tro egen Bull
		-- Robert Burns

%
C, n:Ett programmeringsspråk som är ungefär som Pascal utom mer sommontering förutom att det är inte så mycket som antingen en eller någotannat. Det är antingen det bästa språket tillgängligt för konst idag, ellerdet inte är.
		-- Ray Simard

%
Kål, n .:En välbekant köksträdgård grönsaker ungefär lika stor och klok somen mans huvud.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
cache:En mycket dyr del av minnessystemet för en dator som inte enär tänkt att veta är där.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cahn s Axiom:När allt annat misslyckas, läs instruktionerna.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Campbell lag:Naturen avskyr en innehållslösa försöksledaren.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kanada Bill Jones Motto:Det är moraliskt fel att tillåta rotskott att behålla sina pengar.Kanada Bill Jones Tillägg:En Smith and Wesson slår fyra ess.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Canonical, adj .:Den vanliga eller standard tillstånd eller sätt av något. En sann historia:En Bob Sjöberg, ny på MIT AI Lab, uttryckte några irritation vid användningjargong. Under hans högljudda invändningar, gjorde vi en punkt att använda jargong sommycket som möjligt i sin närvaro, och så småningom började det sjunka in.Slutligen, i en konversation, använde han ordet "canonical" i jargong liknandemode utan att tänka.Steele: "! Aha Vi har slutligen fick du prata jargong för"Stallman: "Vad sa han?"Steele: "Han använde bara 'kanoniska" i den kanoniska sätt. "
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kapten Penny lag:Du kan lura alla människor en del av tiden, ochnågra av de människor hela tiden, men du inte kan lura mamma.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Carperpetuation (kar 'pur husdjur u en shun), n .:Lagen, när du dammsuger, att köra över en sträng åtminstone endussin gånger och nådde över och plocka upp, undersöka det, dåsätta tillbaka ner för att ge vakuum ytterligare en chans.
		-- Rich Hall, "Sniglets"

%
Carsons Tröst:Ingenting är någonsin ett fullständigt misslyckande.Det kan alltid användas som ett dåligt exempel.
		-- Rich Hall, "Sniglets"

%
Carsons Observation på skor:Om skon passar, köpa den andra också.
		-- Rich Hall, "Sniglets"

%
Carswell s Korollarium:När man kommer upp med en bättre råttfälla,natur kommer alltid upp med en bättre mus.
		-- Rich Hall, "Sniglets"

%
Katt, n .:Lapwarmer med inbyggd summer.
		-- Rich Hall, "Sniglets"

%
cerebral atrofi, n:De fenomen som inträffar hjärnceller blir svaga och sjuka, ochförsämra hjärnans prestanda. Ett överflöd av dessa "dåliga" celler kan orsakasymptom relaterade till senilitet, apati, depression och övergripande dålig akademiskaprestanda. Ett visst litet antal hjärnceller kommer att försämras på grund avprestera aktivitet, men stora mängder försvagas av intensiv mental ansträngningoch assimilering av svåra begrepp. Många studenter bliroffer för denna fruktan sjukdom på grund av dåliga vanor såsom overstudying.cerebral darwinism, n:Teorin att effekterna av cerebral atrofi kan vändasgenom renings verkan av tung alkoholkonsumtion. Stora mängder avalkohol orsakar många hjärnceller att dö på grund av syrebrist. Genomprocessen för det naturliga urvalet, kommer de svaga och sjuka hjärnceller dörförsta, bara lämna friska celler. Denna underbara process lämnarimbiber med en friskare, mer levande hjärna, och ökar mental kapacitet.Således är de förödande effekterna av cerebral atrofi vänt och akademiskaprestanda ökar faktiskt bortom tidigare nivåer.
		-- Rich Hall, "Sniglets"

%
Chamberlains lagar:(1) De stora killarna vinner alltid.(2) Allt smakar mer eller mindre som kyckling.
		-- Rich Hall, "Sniglets"

%
teckentäthet, n .:Antalet mycket konstiga människor på kontoret.
		-- Rich Hall, "Sniglets"

%
Välgörenhet, n .:En sak som börjar hemma och oftast stannar där.
		-- Rich Hall, "Sniglets"

%
checkuary, n:Den trettonde månaden på året. Börjar nyårsdagen och slutarnär en person slutar rött skriva det gamla året på sina kontroller.
		-- Rich Hall, "Sniglets"

%
Kock, n .:Någon kock som svär på franska.
		-- Rich Hall, "Sniglets"

%
Cheit klagan:Om du hjälpa en vän i nöd, är han säker på att komma ihåg dig--nästa gång han är i nöd.
		-- Rich Hall, "Sniglets"

%
Kemikalier, n .:Skadliga ämnen från vilka moderna livsmedel görs.
		-- Rich Hall, "Sniglets"

%
Cheops 'lag:Ingenting någonsin blir byggd på schemat eller inom budget.
		-- Rich Hall, "Sniglets"

%
Chicago Transit Authority Rider härskar # 36:Aldrig någonsin be tuffa ser herre bär El Rukn huvudbonaderdär han fick sin "pyramid drivs pizza varmare".
		-- Chicago Reader 3/27/81

%
Chicago Transit Authority Rider härskar # 84:CTA har gratis pop-up timer finns på begäranför överhettade passagerare. När timern dyker upp, förarenglatt baste dig.
		-- Chicago Reader 5/28/82

%
Kycklingsoppa:En gammal mirakelmedicin som innehåller lika delar av AUREOMYCIN,kokain, interferon, och TLC. Den enda krämpa kycklingsoppakan inte bota är neurotiska beroende av en mor.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Chism lag av avslutnings:Den tid som krävs för att slutföra ett statligt projekt ärexakt lika med den tid som redan tillbringat på den.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Chisolm första konsekvens av Murphys andra lag:När saker bara kan omöjligen bli värre, kommer de.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Jul:En dag avskilt av vissa som en tid för kalkon, presenter, tranbärsallader, familj, gemenskap, för andra, noteras som har den bästasvarstiden för hela året.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Churchills Kommentar till Man:Man kommer emellanåt snubblar över sanningen,men för det mesta han kommer att plocka själv upp och fortsätta.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Cinemuck, n .:Kombinationen av popcorn, läsk och smält choklad somtäcker golven i biografer.
		-- Rich Hall, "Sniglets"

%
clairvoyant, n .:En person, vanligtvis en kvinna, som har befogenhet att kontrollera attsom är osynlig för sin beskyddare - nämligen att han är en dumskalle.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Clarkes Slutsats:Låt aldrig din känsla av moral störa göra det rätta.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Clay slutsats:Kreativitet är stor, men plagiat är snabbare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
klon, n:1. En exakt kopia, som i "vår produkt är en klon av derasprodukt. "2. En luddiga, falsk kopia, som i" sin produktär en klon av vår produkt. "
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Clovis "Behandling av en atmosfärisk Anomaly:Den perversa naturen är ingenstans bättre visatän av det faktum att, när den utsätts för samma atmosfär,bröd blir hårt medan kex blir mjuk.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
COBOL:En övning i Artificiell inelegance.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
COBOL:Helt över och bortom förnuftet eller Logic.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cohens lag:Det finns ingen botten till värre.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cohns lag:Ju mer tid du spenderar i rapporteringen om vad du gör, desto mindregång du behöver göra någonting. Stabilitet uppnås när du spenderarall din tid rapportera om ingenting du gör.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kyla, adj .:När politikerna gå omkring med händerna i sina egna fickor.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cole lag:Tunt skivad kål.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Samarbete, n .:En litterär partnerskap som bygger på det felaktiga antagandet attandra kolleger kan stava.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
College:Fontäner av kunskap, där alla går att dricka.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Colvard logiska lokaler:Alla sannolikheter är 50%.Antingen en sak kommer att hända eller det kommer inte.Colvard s unconscionable Kommentar:Detta är särskilt sant när det handlar om någon som du är attraherad av.Grelb s Kommentar:Sannolikheterna är dock 90% mot dig.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Command, n .:Uttalande från en människa och accepterat av en dator iett sådant sätt att den mänskliga känslan som om han är i kontroll.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
kommentar:En överflödig del av det ursprungliga programmet ingår såprogrammerare kan komma ihåg vad fan det var han gjordesex månader senare. Endast den svaga sinnade behöver dem, enligttill dem som tror att de inte är det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Engagemang, n .:[Skillnaden mellan engagemang och] Engagemang kan varaillustreras av en frukost med skinka och ägg. Kycklingen varinblandade, var grisen begåtts.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Utskottet Regler:(1) anländer aldrig på tid, eller du kommer att stämplas en nybörjare.(2) inte säga något förrän mötet är hälften under; dettafrimärken när du är klok.(3) Var så vag som möjligt; detta förhindrar irriterandeandra.(4) Om du är osäker, tyder på att en underkommitté utses.(5) Var först med att flytta för uppskjutande; Detta gör dupopulärt - det är vad alla väntar på.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kommitté, n .:En grupp av män som individuellt kan göra något annat än som en gruppbesluta att ingenting kan göras.
		-- Fred Allen

%
Borgar tre lagar ekologi:(1) Ingen åtgärd är utan biverkningar.(2) Ingenting går någonsin bort.(3) Det finns ingen fri lunch.
		-- Fred Allen

%
Komplext system:En med verkliga problem och imaginära vinster.
		-- Fred Allen

%
Compliment, n .:När du säger något till en annan som alla vet är inte sant.
		-- Fred Allen

%
compuberty, n:Den obekväma period av känslomässiga och hormonella förändringar endator upplevde operativsystemet uppgraderas ochen sun4 sätts delningsfiler.
		-- Fred Allen

%
Datavetenskap:(1) En studie liknar numerologi och astrologi, men saknarprecision av den förra och framgången för den senare.(2) Den utdragna värdeanalys av algoritmer.(3) Den kostsamma uppräkning av det uppenbara.(4) Den tråkiga konsten att hantera ett stort antal trivialiteter.(5) Tautologi utnyttjas i människans tjänst vid ljusets hastighet.(6) The Post-Turing nedgång i formella systemteori.
		-- Fred Allen

%
Dator, n .:En elektronisk enhet som verkställer sekvenser på användbara steg i enhelt förståeligt, noggrant logiskt sätt. Om du trordetta, se mig om en bro jag har till salu på Manhattan.
		-- Fred Allen

%
Koncept, n .:Alla "idé", för vilken en extern konsult faktureras dig mer än$ 25.000.
		-- Fred Allen

%
Konferens, n .:Ett särskilt möte där chefen samlar underlydande att höravad de har att säga, så länge det inte strider mot vadhan redan bestämt sig för att göra.
		-- Fred Allen

%
Förtrogen, förtrogna, n:En anförtros av A med hemligheter B, anför sig genom C.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bekräftat ungkarl:En man som går genom livet utan problem.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Gissningar: Alla udda nummer är prime.Matematiker Bevis:3 är ett primtal. 5 är ett primtal. 7 är ett primtal. Genom induktion, allaudda nummer är prime.Fysiker s Bevis:3 är ett primtal. 5 är ett primtal. 7 är ett primtal. 9 är experimentellfel. 11 är ett primtal. 13 är utmärkt ...Teknikerns Bevis:3 är ett primtal. 5 är ett primtal. 7 är ett primtal. 9 är ett primtal.11 är ett primtal. 13 är utmärkt ...Computer Forskare är ett bevis:3 är ett primtal. 3 är ett primtal. 3 är ett primtal. 3 är prime ...
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Connector Conspiracy, n:[Förmodligen kom in i prominens med utseendet på KL-10,ingen av vars kontakter matchar något annat] Tendensen hostillverkare (eller i förlängningen programmerare eller försäljare av något)att komma med nya produkter som inte passar ihop med den gamlasaker, vilket gör du köper antingen alla nya saker eller dyrtgränssnittsanordningar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Samtycke dekret:Ett dokument där en olycklig företag samtycker att aldrig begåi framtiden oavsett avskyvärda brott mot federal lag detaldrig medgav i första hand.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Konsult, n .:(1) Någon du betalar för att ta klockan från handleden och berättadu vad klockan är. (2) (För återuppta användning) Arbetsnamnetav någon som inte för närvarande innehar ett jobb. Motto: HaKalkylator, Will Travel.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Konsult, n .:[Från con "att bedra, dupera, svindel", eller, möjligen, franska con(Vulgärt) "en person liten förtjänst" + tatet elliptisk form av"Förolämpning."] En tipsaren förklädd som ett orakel, särskilt en somhar lärt sig att decamp vid hög hastighet trots en stor portföljoch tung plånbok.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Konsult, n .:En vanlig människa långt hemifrån.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
konsult, n .:Någon som knowns 101 sätt att älska, men kan inte få ett datum.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Konsult, n .:Någon som hellre klättra i träd och ljuga än att stå påmarken och berätta sanningen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Konsultation, n .:Medicinsk term som betyder "att dela rikedom."
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Konversation, n .:En sång tävling där den som fångar andankallas lyssnaren.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Conway lag:I varje organisation kommer det alltid att finnas en person som vet	vad händer.Denna person måste avfyras.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kopieringsmaskin, n .:En anordning som strimlar papper, blinkar mystiskt kodade meddelanden,och gör dubbletter för alla på kontoret som inteintresserade av att läsa dem.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Corona, n .:Ceremonin att investera en suverän med den yttre och synligatecken på hans gudomliga rätt att blåsas skyhigh med en dynamit bomb.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Korrespondens Korollarium:Ett experiment kan betraktas som en framgång om inte mer än hälftendata måste kasseras för att erhålla korrespondens med din teori.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Corry lag:Papper är alltid starkast vid perforeringarna.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
domstol, n .:En plats där man undvara rättvisa.
		-- Arthur Train

%
Coward, n .:Den som i en farlig akut tänker med benen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Borgenär, n .:En man som har ett bättre minne än en gäldenär.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Crenna lag av politiska ansvar:Om du är den första som får veta om något dåligt, kommer ni att varaansvarig för att agera på det, oavsett din formella arbetsuppgifter.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
kritiker, n .:En person som har själv svårt att tillfredsställa eftersom ingen försökeratt tillfredsställa honom.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Croll s Query:Om tin whistle är gjorda av tenn, vad mistlurar gjord av?
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cropp lag:Mängden arbete varierar inversly med tiden ikontor.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cruickshank lag av kommittéer:Om ett utskott är tillåtet att diskutera en dålig idé tillräckligt länge, detkommer oundvikligen att besluta att genomföra idén helt enkelt eftersom såmycket arbete har redan gjorts på det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
markören adress, n:"Hej, markör!"
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Markör, n .:En vars program kan inte köras.
		-- Robb Russon

%
curtation, n .:Påtvingade komprimering av en sträng i fast längd fältmiljö.Problemet med montering extremt variabel längd strängar såsom namn,adresser, och artikelbeskrivningar i poster med fast längd är ingen trivialmateria. Försummelse av den subtila konsten att curtation har förmodligen fjärmat mermänniskor än någon annan aspekt av databehandling. Du beställer Mozarts "DonGiovanni "från din post klubb, och de fakturera dig $ 24.95 för MOZ DONG.Den witless kartläggning av det sublima till det löjliga! Lika förbryllande ärden curtation som ger samma åtta tecken, det bäst, om duFör "The Best of Wagner", "The Best of Schubert", eller "The Best of the Turds".På samma sätt, vinälskare köper från datoriserade vingårdar snurra sina glasögon,kontrollera sina följesedlar, och informera sina vänner, "En ganska oskyldiga,möjligen overtruncated CAB Sauv 69 TAL. "The klämning av frukten i 10kolumner har gett sådana minnesvärda obsceniteter som COX eller PIP. exemplenciterade är verkliga och curtational metod som producerade dem är fortfarandemed oss.MOZ DONG n.Curtation av Don Giovanni av Wolfgang Amadeus Mozart och Lorenzo daPonte, som utförs av det datoriserade fakturerings ensemble av Internat'lPreview Society, Great Neck (sic), N.Y.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Cutler Webster lag:Det finns två sidor till varje argument, om en personär personligen involverad, i vilket fall det är bara en.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Cyniker, n .:En skurk vars felaktig syn ser saker som de är, intesom de borde vara. Därför anpassade bland skyterna för plockningut en cyniker ögon för att förbättra sin syn.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cyniker, n .:Upplevt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Cyniker, n .:En som ser genom rosafärgade glasögon med en fördomsfull öga.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Data, n .:En periodisering av sugrör på ryggen av teorier.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Data, n .:Computerspeak för "information". korrekt uttalashur Bostonians uttala ordet för ett flickebarn.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Davis lag trafiktäthet:Densiteten för rusningstrafik är direkt proportionell mot1,5 gånger så mycket extra tid du tillåter att komma fram i tid.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Davis Dictum:Problem som försvinner av sig själva, kom tillbaka av sig själva.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Gryning, n .:Den tid då män förnuftets gå till sängs.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Deadwood, n .:Alla i företaget som är mer högre än vad du är.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Death wish, n .:Den enda önskan som alltid går i uppfyllelse, oavsett om man önskar det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Beslutsfattare, n .:Den person på kontoret som var oförmögen att bilda en arbetsgruppinnan musiken stoppas.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
standard N .:[Möjligen från Black engelska "De fel wid DIS systemet är du,vanligare. "] Det fåfängt försök att undvika fel av inaktivitet." Ingenting kommer attkommer ingenting: tala igen "- Kung Lear..
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Standard, n .:Hårdvaran är, naturligtvis.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Deja vu:. Franska, redan sett; inte original; banal.Psychol., Illusionen av att ha tidigare upplevtnågot som faktiskt uppstått för första gången.Psychol., Illusionen av att ha tidigare upplevtnågot som faktiskt uppstått för första gången.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Överläggning, n .:Handlingen att undersöka ett bröd för att avgöra vilken sida det ärsmörade på.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Tandläkare, n .:En JONGLÖR som sätter metall i munnen, drarmynt av sina fickor.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Denver, n .:En ganska liten stad som ligger strax under det så kallade O "i Colorado.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
design, v .:Vad du ångrar inte att göra senare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
DeVries 'dilemma:Om du träffar två knapparna på skrivmaskin, det du inte villträffar papperet.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Dibble första lag Sociologiska:Vissa gör, vissa inte.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Dö, v .:Att sluta synda plötsligt.
		-- Elbert Hubbard

%
Middag förslag # 302 (Hacker De-lite):1 burk importerad skarpsill sardiner i tomatsåsEn påse choklad Malt Carnation Omedelbar frukostEn kartong mjölk
		-- Elbert Hubbard

%
diplomati, n:Ligga i staten.
		-- Elbert Hubbard

%
Dirksen s tre lagarna av politik:(1) bli vald.(2) bli omvald.(3) inte arg, få ännu.
		-- Sen. Everett Dirksen

%
disbar, n:Till skillnad från vissa andra bar.
		-- Sen. Everett Dirksen

%
Distinkt, adj .:En annan färg eller form än våra konkurrenter.
		-- Sen. Everett Dirksen

%
Distress, n .:En sjukdom som uppkommit efter exponering för välstånd en vän.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
skilsmässa, n:En förändring av hustru.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Dokumentation:Instruktioner översatta från svenska från japanska till engelskatalande personer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
dubbelblind experiment, n:Ett experiment där den främsta forskaren tror han ärlurar både motivet och labbassistent. ofta tillsammansav en stark tro på tandfen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Dow lag:I en hierarkisk organisation, ju högre nivå,ju större förvirring.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Drakenberg Discovery:Om du inte tycks kunna hitta dina glasögon,Det är förmodligen för att du inte har dem på.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Drew lag Highway Biology:Det första felet att träffa en ren vindruta landar direkt framfördina ögon.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
drog, n:Ett ämne som, injiceras i en råtta, ger en vetenskaplig uppsats.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ducharme s Precept:Opportunity knackar alltid åtminstone lämpligt tillfälle.Ducharme s Axiom:Om du visar ditt problem tillräckligt nära du kommer att känna igensjälv som en del av problemet.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Tull, n:Vad man förväntar sig från andra.
		-- Oscar Wilde

%
Eagleson lag:Någon kod av din egen att du inte har tittat på för sex eller mermånader, kunde lika gärna ha skrivits av någon annan. (Eaglesonär en optimist, är det verkliga antalet mer som tre veckor.)
		-- Oscar Wilde

%
ekonomi, n .:Ekonomi är läran om värdet och betydelsen av J. K. Galbraith.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Skalfördelar:Uppfattningen att större är bättre. I synnerhet att om du villen viss mängd datorkraft, är det mycket bättre att köpa enbiggie än ett gäng smallies. Accepteras som en trosartikelav människor som älskar stora maskiner och all denna komplexitet. avvisassom en trosartikel av dem som älskar små maskiner och alladessa begränsningar.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
ekonom, n:Någon som är bra med siffror, men har inte tillräckligtpersonlighet för att bli en revisor.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Egotism, n:Gör New York Times korsord med en penna.Egotist, n:En person med låg smak, mer intresserad av sig själv än mig.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ehrman: s kommentar:(1) det kommer att bli värre innan det blir bättre.(2) Vem har sagt det skulle bli bättre?
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Elbonics, n .:De åtgärder på två personer manövrera för ett armstöd i en filmteater.
		-- "Sniglets", Rich Hall & Friends

%
Elchock, n .:Burning på bål med alla moderna förbättringar.
		-- "Sniglets", Rich Hall & Friends

%
Elefant, n .:En mus byggd för statliga specifikationer.
		-- "Sniglets", Rich Hall & Friends

%
Elfte lag akustik:I en minsta-fassystem det finns ett oupplösligt samband mellanfrekvensomfång, fas respons och övergående svar, eftersom deär alla bara förvandlas av varandra. Detta i kombination medminimalization av öppen slinga fel i utgångsförstärkare och korrektersättning för icke-linjära passiva delningsfilter belastning kanleda till en betydande minskning av systemets upplösning förlorad. Dock,naturligtvis allt detta betyder uttaget när du lyssnar på Pink Floyd.
		-- "Sniglets", Rich Hall & Friends

%
Emacs, n .:En långsam parodi av en textredigerare.
		-- "Sniglets", Rich Hall & Friends

%
Emersons lag motsatsförhållande:Vår främsta vill i livet är någon som ska få oss att göra vad vikan. Ha funnit dem, ska vi då hatar dem för det.
		-- "Sniglets", Rich Hall & Friends

%
Encyclopedia Salesmen:Bjuda in dem alla i. Kväva ut bakvägen. Ring polisenoch berätta ditt hus är inbrott.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Ändlös slinga, n .:se Loop, Endless.Loop, Endless, n .:se oändlig loop.
		-- Random Shack Data Processing Dictionary

%
Engram, n .:1. Den fysiska manifestationen av människans minne - "engrammet."2. En särskild minne i fysisk form. [Användning anmärkning: denna term är inte längrei allmänt bruk. Före Wilson och Magruder historiska upptäckt, naturenav engrammet var ett ämne för intensiv spekulation bland neuroforskare,psykologer och även datavetare. 1994 Professorer M. R. Wilsonoch W. V. Magruder båda Mount St Coax University i Palo Alto, visadeslutgiltigt att däggdjurshjärnan är hårdkodade att tolka en uppsättningtrettio sju genetiskt överförda samarbetsvilliga TECO makron. mänskliga minnetvisade att uppehålla sig i 1 miljon Q-register som Huffman kodad enbart versalerASCII-strängar. Intresset för engram har minskat väsentligt sedan desstid.]3: e upplagan, 2007 A.D.
		-- New Century Unabridged English Dictionary,

%
förbättra, v .:Att manipulera en bild, vanligen till skada.
		-- New Century Unabridged English Dictionary,

%
Entreprenuer, n .:En hög-rullande risktagare som hellrevara ett spektakulärt misslyckande än en dyster framgång.
		-- New Century Unabridged English Dictionary,

%
Avund, n .:Önskar du hade fötts med en orättvis fördel,istället för att behöva försöka förvärva en.
		-- New Century Unabridged English Dictionary,

%
Epperson lag:När en man säger att det är en dum, barnslig lek, det är nognågot som hans hustru kan slå honom på.
		-- New Century Unabridged English Dictionary,

%
Etymologi, n .:Några tidiga etymologiska forskare kom upp med avledningar somvar svårt för allmänheten att tro. Uttrycket "etymologi" bildadesfrån latinets "etus" ( "ätit"), roten "mal" ( "dåligt"), och "nik"	("studie av"). Det betydde "studiet av saker som är svåra att svälja."
		-- Mike Kellen

%
Varje häst har ett oändligt antal ben (bevis genom hotelser):Hästar har ett jämnt antal ben. Bakom de har två ben, och ifront de har fore-ben. Detta gör sex ben, som visserligen är enudda antal ben för en häst. Men det enda numret som är både medoch udda är oändligheten. Därför hästar har ett oändligt antalben. Nu för att visa detta för det allmänna fallet anta att någonstans,det finns en häst som har ett ändligt antal ben. Men det är en hästav annan färg, och lemmat [ "Alla hästar har samma färg"]som inte existerar.
		-- Mike Kellen

%
Varje program har (minst) två syften:den för vilken den skrevs och en annan som inte var det.
		-- Mike Kellen

%
Bekostnad konton, n .:Corporate matkuponger.
		-- Mike Kellen

%
Erfarenhet, n .:Något du inte får förrän strax efter att du behöver det.
		-- Olivier

%
Expert, N .:Någon som kommer ut ur staden och visar bilder.
		-- Olivier

%
Utdrag från Official Utlottning Regler:INGEN köp krävs för att få din PRISAtt göra anspråk på din vinst utan inköp, gör följande: (a) försiktigtklippa ut datorn tryckt namn och adress från övre högrahörnet av priset kravformuläret. (B) Montera datornamnförtydligande ochadress - med lim eller tejp (inga häftklamrar eller gem) -till en 3x5 tum indexkort. (C) snitt också in "Nej" punkt (lägrevänstra hörnet av Prize krav Form) och fäst den på 3x5 kortunder din adressetikett. (D) därefter ut på 3x5 kort, ovanfördator tryckta namn och adress orden "CARTER & VAN PEELSWEEPSTAKE "(Använd stora bokstäver.) (E) Slutligen placera 3x5 kort(Utan att böja) i en vanlig kuvert [OBS: använd inte det denOfficiell Prize krav och CVP Parfym svarskuvert eller så kan du varadiskvalificerad], och post till: CVP, Box 1320, Westbury, NY 11595. Skriv utden här adressen korrekt. Följa ovanstående instruktioner noga ochhelt eller så kan du diskvalificeras från att ta emot ditt pris.
		-- Olivier

%
Saga, n .:En skräckhistoria att förbereda barnen för tidningarna.
		-- Olivier

%
Fakir, n:En psykolog vars karismatiska uppgifter har inspirerat nästanreligiös hängivenhet i hans anhängare, även om källornaverkar ha shinnied upp ett rep och försvann.
		-- Olivier

%
falsie försäljare, n:Fylligare byst man.
		-- Olivier

%
Kända sista ord:
		-- Olivier

%
Kända sista ord:(1) "Oroa dig inte, jag klarar det."(2) "Du och vilken armé?"(3) "Om du var lika smart som du tror att du är, du skulle inte varaen polis. "
		-- Olivier

%
Kända sista ord:(1) Dra inte ut det, kommer det bara ta en stund att åtgärda.(2) Låt oss ta en genväg, kan han inte se oss därifrån.(3) Vad händer om du rör dessa två trådar tog--(4) Vi kommer inte behöver reservationer.(5) Det är alltid soligt det den här tiden på året.(6) Oroa dig inte, det är inte laddad.(7) De skulle aldrig (vara dum nog att) göra honom en chef.(8) inte orolig! Kvinnor älskar det!
		-- Olivier

%
Kända citat:""""""
		-- Marcel Marceau

%
Kända, adj .:Iögonfallande olycklig.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
funktionen, n:En överraskande egenskap hos ett program. Occasionaly dokumenteras. Tillkalla en fastighet en funktion innebär ibland författaren inteöverväga det fallet, och programmet gör en oväntad, meninte nödvändigtvis fel svar. Se BUG. "Det är inte en bugg, det ären funktion! "En bugg kan ändras till en funktion genom att dokumentera den.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
fenderberg, n .:De stora glaciala avlagringar som bildas på insidanöver bil fendrar under snöstormar.
		-- "Sniglets", Rich Hall & Friends

%
Fergusons Precept:En kris är när du inte kan säga "låt oss glömma alltihop."
		-- "Sniglets", Rich Hall & Friends

%
Fidelity, n .:En förtjänst är utmärkande för dem som är på väg att bli förrådd.
		-- "Sniglets", Rich Hall & Friends

%
Femte lag tillämpad Terror:Om du får en öppen bok examen, kommer du att glömma din bok.Naturlig följd:Om du får en hemtentamen, kommer du att glömma var du bor.
		-- "Sniglets", Rich Hall & Friends

%
Femte lag förhalning:Förhalning undviker ledan; en har aldrig en känsla av attdet finns inget viktigt att göra.
		-- "Sniglets", Rich Hall & Friends

%
Arkivskåp:En fyra låda, aktiveras manuellt papperskorgen komprimator.
		-- "Sniglets", Rich Hall & Friends

%
filibuster, n .:Kasta din vänta.
		-- "Sniglets", Rich Hall & Friends

%
Finagle s Creed:Vetenskap är sant. Inte vilseledas av fakta.
		-- "Sniglets", Rich Hall & Friends

%
Finagle åttonde lag:Om ett experiment fungerar har något gått fel.Finagle nionde lag:Oavsett vad resultat förväntas, är alltid beredda att någon	låtsas.Finagle tionde lag:Oavsett vad resultatet någon är alltid angelägna om att misstolka det.Finagle elfte lag:Oavsett vad som händer, tror någon det hände enligthans husdjur teori.
		-- "Sniglets", Rich Hall & Friends

%
Finagle första lag:Om ett experiment fungerar har något gått fel.
		-- "Sniglets", Rich Hall & Friends

%
Finagle första lag:För att studera ett ämne bäst förstår det ordentligt innan du börjar.Finagle andra lag:alltid hålla ett register över uppgifter - det visar att du har arbetat.Finagle fjärde lag:När ett jobb sotigt upp, något göras för att förbättra det bara gördet värre.Finagle femte lag:Dra alltid dina kurvor, sedan rita dina avläsningar.Finagle sjätte lag:Tror inte på mirakel - lita på dem.
		-- "Sniglets", Rich Hall & Friends

%
Finagle andra lag:Oavsett vad den förväntade resultat, kommer det alltid att finnasnågon ivrig att (a) misstolka den, (b) fejka det, eller (c) anser att dethände enligt hans eget husdjur teori.
		-- "Sniglets", Rich Hall & Friends

%
Finagle sjunde lag:Den perversa universum tenderar mot ett maximum.
		-- "Sniglets", Rich Hall & Friends

%
Finagle tredje lag:I varje insamling av uppgifter, siffran mest uppenbart rätt,bortom allt behov av kontroll, är misstagetkorollarier:(1) Ingen vem du ber om hjälp kommer att se det.(2) Den första personen som stannar, vars råd du verkligeninte vill höra, kommer att se det omedelbart.
		-- "Sniglets", Rich Hall & Friends

%
Fina s Korollarium:Funktionalitet föder förakt.
		-- "Sniglets", Rich Hall & Friends

%
Finster lag:En stängd mun samlar ingen fot.
		-- "Sniglets", Rich Hall & Friends

%
Första lag Cykel:Oavsett vilken väg du rida, det är uppförsbacke och motvind.
		-- "Sniglets", Rich Hall & Friends

%
Första lag debatt:Aldrig argumentera med en idiot. Folk kanske inte vet skillnaden.
		-- "Sniglets", Rich Hall & Friends

%
Första lag förhalning:Förhalning förkortar jobbet och lägger ansvaretför sin uppsägning på någon annan (dvs. den myndighet sominförde tidsfristen).Femte lag förhalning:Förhalning undviker ledan; en har aldrig en känsla av attdet finns inget viktigt att göra.
		-- "Sniglets", Rich Hall & Friends

%
Första lag socio Genetics:Celibat är inte ärftlig.
		-- "Sniglets", Rich Hall & Friends

%
Första Rule of History:Historia upprepar sig inte - historiker bara upprepa varandra.
		-- "Sniglets", Rich Hall & Friends

%
Fiskskål, n .:En inglasade isoleringscell där nyligen främjas cheferhålls för observation.
		-- "Sniglets", Rich Hall & Friends

%
Fem regler för evigt elände:(1) Försök alltid att uppmana andra att titta på dig positivt.(2) Gör massor av antaganden om situationer och se till attbehandla dessa antaganden som om de är verklighet.(3) Sedan behandla varje ny situation som om det är en kris.(4) leva i det förflutna och bara framtiden (blir besatthur mycket bättre saker kan ha varit eller hur mycket sämresaker kan bli).(5) Ibland stampa på dig själv för att vara så dum attFölj de fyra första regler.
		-- "Sniglets", Rich Hall & Friends

%
flannister, n .:Plast ok som har en sex-pack öl tillsammans.
		-- "Sniglets", Rich Hall & Friends

%
Flon lag:Det finns inte nu, och kommer aldrig att bli, ett språksom är det minsta svårt att skriva dåliga program.
		-- "Sniglets", Rich Hall & Friends

%
flödesschema, n. & V .:[Från flöde "till krusning i rika överflöd, som hår" + kart"Ett kryptiskt dolda skattkarta som syftar till att vilseleda den oinvigde."]1. n. Lösningen, om någon, till en klass av Mascheroni konstruktionproblem där givna algoritmer kräver geometrisk representationmed endast 35 grundläggande ideogram av ANSI mallen. 2. n. Neronicdoodling medan systemet brinner. 3. n. En låg kostnad substitut förtapet. 4. n. Den innumerate vilseledande analfabeter. "ENtusen bilder är värt tio rader kod. "- programmerarensLittle Red vademecum, Mao Tse T'umps. 5. v.intrans. Att produceraflödesscheman utan särskilt syfte i åtanke. 6. v.trans. att fördunkla(Ett problem) med esoteriska karikatyrerna.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Flugg lag:När du behöver ta i trä är när du inseratt världen består av vinyl, Naugahyde och aluminium.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Dimljus, n .:Alltför (ofta obnoxiously) ljusa lampor monterade på fronternaav bilar; användas på torra, klara nätter för att indikera attförarens hjärna är i en dimma. Se även "Idiot Lights".
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Idiotsäker Operation:Ingen avsättning för justering.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Prognos, n .:En förutsägelse om framtiden, baserat på det förflutna, försom prognosmakare kräver betalning i nuet.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Glömska, n .:En gåva från Gud skänkte gäldenärer i kompensation förderas armod av samvete.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
FORTUNE förklarar vad JOBB ÖVERSIKT slagord MEAN: # 1skicklig oral kommunikatör:Mumbles ohörbart när du försöker att tala. Pratar med själv.Argumenterar med själv. Förlorar dessa argument.skicklig skriven kommunikatör:Klotter väl. Teckningar är oföränderliga oläsliga, med undantag förde delar som tillskriver de senaste misslyckanden till någon annan.tillväxtpotential:Med rätt vägledning, återkommande rådgivning och stödundervisning,den reviewee kan ges tillräckligt med tid och noggrann övervakning, träffade minimikrav som förväntas av honom från bolagets sida.nyckel företag siffra:Fungerar som den perfekta motexempel.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
FORTUNE förklarar vad JOBB ÖVERSIKT slagord MEAN: # 4konsekvent:Reviewee har inte fått något rätt ännu, och det förväntasatt detta mönster kommer att fortsätta under det kommande året.en utmärkt bollplank:Nuvarande reviewee med valfritt antal alternativ, och genomföradem i den ordning precis motsatsen till hans / hennes specifikation.en planerare och organisatör:Vanligtvis lyckas sätta på strumpor innan skor. Kan matchadjur taggar på hans kläder.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
FORTUNE förklarar vad JOBB ÖVERSIKT slagord MEAN: # 9har ledningen potential:På grund av hans intima relation med döda ting, denreviewee har utsetts till den kritiska läget för avdelningenpenna monitor.inspirerande:En sann inspiration för andra. ( "Där men för Guds nåd,gå I. ")anpassar sig till stress:Passerar vind, vatten, eller ut beroende på svårighetsgraden avsituation.målinriktad:Ständigt sätter låga mål för sig själv, och oftast misslyckasatt möta dem.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Fortune Regler för Memo Wars: # 2Med tanke på de otroliga framsteg inom sociocybernetics och telepsychology överde senaste åren, kan vi nu att helt förstå allt somförfattaren av en PM försöker säga. Tack vare moderna utvecklingeni electrocommunications som anteckningar, vnews och el, har vi enotrolig nivå av interunderstanding vars like civilisationen haraldrig känt. Således, annars finns risk för att din misstolka någonmemo är praktiskt taget noll. Att veta detta, någon som anklagar dig för att hagjort så är en lögnare, och bör behandlas därefter. Om du * gör * förståPM i fråga, men har absolut ingenting av substans att säga,du har ett utmärkt tillfälle för en ond ad hominem attack. Faktiskt,de enda * olämpliga * gånger för en ad hominem attack är som följer:1: När du håller helt med författaren av en PM.2: När författaren av den ursprungliga PM är mycket större än vad du är.3: När du svarar på en av dina egna anteckningar.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Fjärde lag tillämpad Terror:Natten innan engelsk historia halvtids din biologiinstruktör kommer att tilldela 200 sidor om planaria.Naturlig följd:Varje instruktör förutsätter att du har ingenting annat att göra än attstudera för att instruktörskurs.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Fjärde lag Revision:Det är oftast opraktiskt att oroa i förväg omstörningar - om du har någon, kommer någon att göra något för dig.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Fjärde termodynamikens:Om sannolikheten för framgång är inte nästan ett, är det fan nära noll.
		-- David Ellis

%
Fresco Discovery:Om du visste vad du gjorde skulle du förmodligen vara uttråkad.
		-- David Ellis

%
Fried 1st regel:Ökad automatisering av kontorsarbete funktionalltid leder till ökade driftskostnader.
		-- David Ellis

%
Vänner, n .:Folk som lånar dina böcker och som våta glasögon på dem.Personer som känner dig väl, men gillar dig ändå.
		-- David Ellis

%
Frobnicate, v .:Att manipulera eller justera för att justera. Härstammar från FROBNITZ. Vanligtvisförkortat till FROB. Således en har talesättet "att FROB en FROB." se TWEAKoch twiddle. Användning: FROB, rulla och justera ibland beteckna punkter längsett kontinuum. FROB connotes aimless manipulation; KRUMELUR connotes bruttomanipulation, ofta en grov sökning för en ordentlig inställning; justera betecknarfinjustering. Om någon vänder en ratt på ett oscilloskop, så om han ärnoggrant anpassa den han förmodligen tweaking det; om han bara vänder detmen titta på skärmen han är nog tråkigt det; men om han är baragör det eftersom att vrida en ratt är roligt, han frobbing det.
		-- David Ellis

%
Frobnitz, pl. Frobnitzem (frob'nitsm) N .:En ospecificerad fysiskt objekt, en widget. hänvisar också till elektroniskasvarta lådor. Denna sällsynt form är vanligtvis förkortat till Frotz, eller mervanligen till FROB. Även använda är FROBNULE, FROBULE och FROBNODULE.Från och kanske 1979, FROBBOZ (Fruh-bahz), pl. FROBBOTZIM, har ocksåblivit mycket populärt, främst på grund av sin exponering via Adventure spin-offkallas Zork (Dungeon). Dessa kan också tillämpas på icke-fysiska föremål,såsom datastrukturer.
		-- David Ellis

%
Fuchs Varning:Om du verkligen ser ut som din passfoto, du är inte branog att resa.
		-- David Ellis

%
Fudd första lag Opposition:Tryck något tillräckligt hårt och det kommer att falla över.
		-- David Ellis

%
Roliga experiment:Få en burk raklödder, kasta den i en frys för ungefär en vecka.Ta sedan ut, dra metallen och sätta den där du vill ...sovrum, bil, etc. Som det tinar, expanderar det en otrolig mängd.
		-- David Ellis

%
Roliga fakta, # 14:I bordtennis, vem får 21 poäng första vinner. Det är hurdet en gång var i baseball - vem fick 21 körningar först vann.
		-- David Ellis

%
Roliga fakta, # 63:Namnet Kalifornien gavs till staten av spanska conquistadorerna.Det var namnet på en imaginär ö, ett paradis på jorden, iSpanska roman "Les Serges de Esplandian", skriven av Montalvo i1510.
		-- David Ellis

%
furbling, v .:Att behöva vandra genom en labyrint av rep på en flygplats eller bankäven när du är den enda personen i linje.
		-- Rich Hall, "Sniglets"

%
Galbraith lag av den mänskliga naturen:Inför valet mellan att ändra sitt sinne och bevisa attfinns det ingen anledning att göra det, blir nästan alla upptagen på bevis.
		-- Rich Hall, "Sniglets"

%
Genderplex, n .:Situationen för en person i en restaurang som är oförmögen attfastställa hans eller hennes utsedda toaletten (t.ex. sköldpaddor).
		-- Rich Hall, "Sniglets"

%
släktforskning, n .:En redogörelse för en härstamning från en förfadersom inte särskilt noga med att spåra sin egen.
		-- Ambrose Bierce

%
Geni, n .:En kemist som upptäcker en tvätttillsats som rimmar med "ljus".
		-- Ambrose Bierce

%
geni, n .:Person smart nog att födas på rätt plats vid rätttidpunkten för rätt kön och att följa upp denna fördel genom att sägaalla de rätta sakerna för alla rätt personer.
		-- Ambrose Bierce

%
genlock, n .:Varför han stannar i flaskan.
		-- Ambrose Bierce

%
Gerrold lagar av Infernal Dynamics:(1) Ett objekt i rörelse kommer alltid att ledas i fel riktning.(2) Ett föremål i vila kommer alltid att vara på fel plats.(3) Den energi som krävs för att ändra antingen en av dessa tillståndkommer alltid att vara mer än du vill förbruka, men aldrig såmycket som för att göra arbetet helt omöjligt.
		-- Ambrose Bierce

%
Få jobbet gjort är ingen ursäkt för att inte följa reglerna.Naturlig följd:Följa reglerna inte kommer att få jobbet gjort.
		-- Ambrose Bierce

%
Gilberts Discovery:Varje försök att använda de nya super lim resulterar i de två delarnaklibba till tummen och pekfingret i stället för till varandra.
		-- Ambrose Bierce

%
Ginsbergs Sats:(1) Du kan inte vinna.(2) Du kan inte nollresultat.(3) Du kan inte ens avsluta spelet.Freemans kommentar på Ginsberg sats:Varje större filosofi som försöker göra livet verkarmeningsfull bygger på negationen av en del av GinsbergsSats. Nämligen:(1) Kapitalismen baseras på antagandet att man kan vinna.(2) Socialismen är baserad på antagandet att du kan gå jämnt ut.(3) Mysticism är baserad på antagandet att man kan avsluta spelet.
		-- Ambrose Bierce

%
Ginsburg lag:I samma ögonblick du tar bort din sko i en skoaffär, dinstortån kommer att dyka ut ur strumpan för att se vad som händer.
		-- Ambrose Bierce

%
gleemites, n .:Förstenade fyndigheter av tandkräm som finns i sänkor.
		-- "Sniglets", Rich Hall & Friends

%
Glib fjärde lag Otillförlitligt:Investeringar i tillförlitlighet kommer att öka tills den överstigertroliga kostnaden för fel, eller tills någon insisterar på att fånågra nyttigt arbete.
		-- "Sniglets", Rich Hall & Friends

%
Gnagloot, n .:En person som lämnar alla sina liftkort på kavajen baraimponera på folk.
		-- Rich Hall, "Sniglets"

%
Goda s Truism:Med den tid du kommer till den punkt där du kan gå ihop,någon flyttar ändarna.
		-- Rich Hall, "Sniglets"

%
Godwins lag (prov [Usenet].):Som en Usenet diskussion blir längre, sannolikheten för enjämförelse involverar nazister eller Hitler närmar en. "Det finns entradition i många grupper som, när detta inträffar, är att trådenöver, och den som nämns nazisterna har automatiskt förloratoavsett argument pågick. Godwins lag garanterar därmedatt det föreligger en övre gräns för gänglängden i dessa grupper.
		-- Rich Hall, "Sniglets"

%
Guld lag:Om skon passar, det är fult.
		-- Rich Hall, "Sniglets"

%
Guld, n .:En mjuk formbar metall relativt sällsynta i distributionen. Detbryts djupt i jorden fattiga män som sedan ge det till rikamän som omedelbart begrava tillbaka i jorden i stora fängelser,även om guld har inte gjort något för dem.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Goldenstern regler:(1) hyra alltid en rik advokat(2) Aldrig köpa från en rik försäljare.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Gomme s lagar:(1) En backscratcher kommer alltid att hitta nya kliar.(2) Tiden accelererar.(3) Vädret hemma förbättras så snart du går bort.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Gordons första lag:Om ett forskningsprojekt är inte värt att göra, är det inte värt att göra väl.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Gordons lag:Om du tror att du har lösningen, var frågan dåligt formulerade.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
skvaller, n .:Höra något du tycker om någon du inte.
		-- Earl Wilson

%
Goto, n .:Ett programmeringsverktyg som finns för att tillåta strukturerade programmerareatt klaga ostrukturerade programmerare.
		-- Ray Simard

%
Regeringens lag:Det finns ett undantag till alla lagar.
		-- Ray Simard

%
Grabel lag:2 inte är lika med tre - inte ens för stora värden på två.
		-- Ray Simard

%
Morfar Charnock lag:Du aldrig riktigt lära sig att svära tills du lära dig att köra.[Jag trodde det var när barnen lärde sig att köra. Ed.]
		-- Ray Simard

%
grasshopotomaus:En varelse som kan hoppa till enorma höjder ... en gång.
		-- Ray Simard

%
Allvar:Vad du får när du äter för mycket och för snabbt.
		-- Ray Simard

%
Gray lag av programmering:`_ N + 1 'triviala uppgifter förväntas ske i sammatid som `_ n 'uppgifter.Logga in på Rebuttal Gray lag:`_ N + 1 'triviala uppgifter tar dubbelt så lång tid som` _ n' triviala uppgifter.
		-- Ray Simard

%
Stor amerikansk Axiom:Vissa är bra, mer är bättre, för mycket är precis lagom.
		-- Ray Simard

%
Greens lag Debatt:Allt är möjligt om du inte vet vad du pratar om.
		-- Ray Simard

%
Greener lag:Aldrig argumentera med en man som köper bläck genom pipan.
		-- Ray Simard

%
Grelb påminnelse:Åttio procent av alla människor anser sig vara ovangenomsnittliga förare.
		-- Ray Simard

%
Griffin tanke:När du svälta med en tiger, svälter tigern sist.
		-- Ray Simard

%
Grinnell lag of Labor slapphet:I alla tider, för alla uppgifter, du har inte fått tillräckligt görs idag.
		-- Ray Simard

%
Giljotin, n .:En fransk hack centrum.
		-- Ray Simard

%
Gumperson lag:Sannolikheten för att en viss händelse inträffar är omväntproportionell mot dess önskvärdhet.
		-- Ray Simard

%
Gunter s Airborne Upptäckter:(1) När du serveras en måltid ombord på ett flygplan,flygplanet kommer att stöta turbulens.(2) Styrkan hos turbulensenär direkt proportionell mot temperaturen i ditt kaffe.
		-- Ray Simard

%
gurmlish, n .:Den röda varningsflagga på toppen av en club sandwich somhindrar personen från att bita i det och punktera taketfrån hans mun.
		-- Rich Hall, "Sniglets"

%
guru, n .:En person i T-shirt och sandaler som tog en hiss rida meden senior vice president och är ytterst ansvarig förtelefonsamtal du är på väg att få från din chef.
		-- Rich Hall, "Sniglets"

%
guru, n:En dator ägare som kan läsa manualen.
		-- Rich Hall, "Sniglets"

%
gyroskop, n .:Ett hjul eller skiva monterad för att snurra snabbt omkring en axel och ävenfri att rotera kring en eller båda av två axlar perpindicular tillvarandra och axeln för dragning, så att en rotation av ett av detvå inbördes vinkelräta axlar resultat från tillämpning avvridmoment till den andra när hjulet snurrar och så attHela apparaten erbjuder betydande motstånd beroende pårörelsemängdsmomentet för alla moment som skulle ändra riktningför axeln för dragning.
		-- Webster's Seventh New Collegiate Dictionary

%
H.L. Mencken lag:De som kan - göra.De som inte kan - undervisa.Martins Extension:De som inte kan lära - Administrera.
		-- Webster's Seventh New Collegiate Dictionary

%
Hacker lag:Tron att ökad förståelse nödvändigtvis rören nation till handling är en av mänsklighetens äldsta illusioner.
		-- Webster's Seventh New Collegiate Dictionary

%
Hacker Quicky # 313:Gräddfil -n- Onion chipsMikrovågsugn Egg Roll	Chokladmjölk
		-- Webster's Seventh New Collegiate Dictionary

%
hacker, n .:En mästare Byter.
		-- Webster's Seventh New Collegiate Dictionary

%
hacker, n .:Ursprungligen varje person med en knack för tvinga envis livlösa	saker; därmed en person med ett lyckligt knack senare kontrakterats av denmytiska filosof Frisbee Frobenius den gemensamma användning, "hacka".I gamla tider, efter slutförandet av vissa särskilt avskyvärda kroppav kodning som hände för att fungera bra, skulle culpable programmerare samlai en liten cirkel runt en första upplagan av Knuth bästa Volym I avlevande ljus, och fortsätt att få mycket berusade medan sporadiskt skärandeföljande sång:Hacker slagsmål SongHan är en Hack! Han är en Hack!Han är en kille med den lyckliga knep!Aldrig förfuskar, aldrig försummar,Alltid blir hans saker att fungera!Alla tar en drink (viktigt!)
		-- Webster's Seventh New Collegiate Dictionary

%
Hale Mail regel:När du är redo att svara på ett brev, kommer du saknar åtminstoneen av följande:(A) En penna eller skrivmaskin.(B) brevpapper.(C) Frimärke.(D) brevet du svarar.
		-- Webster's Seventh New Collegiate Dictionary

%
halv-done, n .:Detta är det bästa sättet att äta en kosher dill - när det är fortfarande krispigt,ljusgrön, men full av vitlök smak. Skillnaden mellan dettaoch den typiska fuktig mörkgrön gurka lik är somskillnaden mellan liv och död.Du kan finna det svårt att hitta en bra halv-done kosher dill däri Seattle, så vad du bör göra är att ta en taxi ut till flygplatsen,flyga till New York, ta JFK Express till Jay Street-Borough Hall,överföra till en uptown F, gå av vid East Broadway, gå norrut påEssex (längs parken), gör din första vänster in på Hester Street, promenadcirka femton steg, vrid nittio grader åt vänster, och stopp. Säg tillman, "Låt mig få en trevlig halv-done." Värt besväret, var inte det?
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Sidan, n .:En singulär instrument bärs vid slutet av en mänsklig arm ochvanligen kastas in någons ficka.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
handskakningsprotokoll, n:En process som används av fientliga externa enheter initiera enbryskt men medborgardialog, vilket i sin tur kännetecknas avenstaka missförstånd, tjura, och utskällningar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Baksmälla, n .:Bevisbördan.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
baksmälla, n .:Vrede av druvor.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hanlon rakkniv:attribut aldrig malice det som adekvat förklarasav stupidity.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hansons Behandling av tid:Det finns aldrig tillräckligt med timmar på en dag, men alltid alltför många dagarinnan lördag.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Lycka, n .:En angenäm känsla som uppstår från överväger elände annan.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
hårt, adj .:Kvaliteten på din egen data; också hur det är att tro demandra människor.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hårdvara, n .:De delar av ett datorsystem som kan sparkas.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Harriets Dining Observation:På varje restaurang, hårdheten hos smör klapparökar i direkt proportion till mjukheten hos brödet.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Harris Lament:Alla de goda tas.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Harrisberger fjärde lag Lab:Erfarenhet är direkt proportionell mot mängden utrustning som förstörd.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Harrison postulatet:För varje handling finns en likvärdig och motsatt kritik.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hartley första lag:Du kan leda en häst till vatten, men om du kan få honom att flytapå ryggen, har du fått något.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hat, n .:En känsla lämpligt att i samband med en annan överlägsenhet.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hawkeye slutsats:Det är inte lätt att spela clown när du har att köra helacirkus.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Himmel, n .:En plats där de ogudaktiga längre från bekymrar dig med tal omderas personliga angelägenheter, och bra lyssna med uppmärksamhet när duförklara din egen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
tung, adj .:Förföras av choklad sidan av kraften.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Heller lag:Den första myten om ledningen är att det existerar.Johnsons Korollarium:Ingen vet riktigt vad som händer var som helst inomorganisation.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hempstone Fråga:Om du måste resa på Titanic, varför inte gå första klass?
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Herth lag:Han som vänder andra kinden för långt blir det i nacken.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hewett Observations:Elakhet av en byråkrat är omvänt proportionell mot hans ellersin ställning i regeringshierarkin och antaletkamrater liknande ingrepp.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hildebrant princip:Om du inte vet vart du ska, kommer alla vägar dit du.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hippogriff, n .:Ett djur (numera utdöd) som var till hälften häst och hälften grip.Gripen var själv en förening varelse, hälften lejon och hälften örn.Hippogriffen var faktiskt därför endast en fjärdedel örn, vilketär två dollar och femtio cent i guld. Studiet av zoologi är fullav överraskningar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Historia, n .:Papa Hegel han säger att allt vi lär av historien är att vilära ingenting av historien. Jag känner folk som inte ens kan lära avvad som hände i morse. Hegel måste ha tagit ett längre perspektiv.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Hitchcocks Staple Princip:Häftapparaten tar slut häftklamrar bara när du försökerstapel något.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Hlade lag:Om du har en svår uppgift, ge det till en lat människa -de kommer att hitta ett enklare sätt att göra det.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Hoare lag av stora problem:Inuti varje stort problem är ett litet problem som kämpar för att komma ut.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Hoffer s Discovery:Den stora handling av en döende institution är att utfärda ett nyttrevideras förstorad upplaga av riktlinjer och rutiner manual.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Hofstadter lag:Det tar alltid längre tid än förväntat, även när du tarHofstadter lag i beräkningen.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Hollerith, v .:Vad du giver när din telefon är på fritzeth.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
smekmånad, n .:En kort period av doting mellan dating och debting.
		-- Ray C. Bandy

%
Honorable, adj .:Lider av ett hinder i en räckhåll. i lagstiftningsorgan, är det brukligt att tala om alla medlemmar som hederlig; som,"Den ärade gentlemannen är en skörbjugg byracka."
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Horners Fem Thumb Postulat:Erfarenheterna varierar direkt med utrustning förstörd.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Horngren Observations:Bland ekonomer, är den verkliga världen ofta ett specialfall.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hushålls tips:Om du är ute ur grädde för ditt kaffe, gör majonnäs endandy substitut.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
HUR DU kan säga att det kommer att bli kärvt:# 1040 inkomst check studsar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
HUR DU kan säga att det kommer att bli kärvt:# 15 Ditt husdjur sten snäpper på dig.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
HUR DU kan säga att det kommer att bli kärvt:# 32: Du kallar din telefonsvarare och de har aldrig hört talas om dig.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Howe lag:Alla har ett system som inte kommer att fungera.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hubbard lag:Ta inte livet för allvarligt; du kommer inte att få ut av det levande.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Hurewitz Memory Princip:Chansen att glömma något är direkt proportionelltill ... till ... eh .....
		-- Ambrose Bierce, "The Devil's Dictionary"

%
IBM Pollyanna Princip:Maskiner ska fungera. Folk borde tänka.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
IBM: s ursprungliga motto:Cogito ergo vendo; Vendo ergo sum.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
IBM:[International Business Machines Corp.] Även känd som Itty BittyMaskiner eller Advokaten vän. Den dominerande kraften i datornmarknadsföring och har levererat över hela världen cirka 75% av alla kända hårdvaraoch 10% av alla program. För att skydda sig från litigious avundmindre framgångsrika organisationer, såsom den amerikanska regeringen, IBMsysselsätter 68% av alla kända ex-advokat Allmänt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
IBM:Jag har flyttatsIdioter bli cheferIdioter Köp merOmöjligt att köpa MachineOtroligt stor maskinBranschens största misstagInternational Brotherhood of MercenariesDet svindlarDet är bättre manuelltItty-Bitty Machines
		-- Ambrose Bierce, "The Devil's Dictionary"

%
IBM:Det kan vara långsam, men det är svårt att använda.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
idiot box, n .:Den del av höljet som berättar en person, om att placerastämpla när de inte riktigt kan lista ut det själva.
		-- Rich Hall, "Sniglets"

%
Idiot, n .:En medlem av en stor och kraftfull stam vars inflytande i människorsfrågor har alltid varit dominerande och kontrollerande.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
sysslolöshet, n .:Fritid gått till utsäde.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
ignisecond, n:Den överlappande tidsögonblick när handen låsa bilendörr även när hjärnan säger, "mina nycklar är där!"
		-- Rich Hall, "Sniglets"

%
okunnighet, n .:När du inte vet någonting, och någon annan får reda på.
		-- Rich Hall, "Sniglets"

%
Iles lag:Det finns alltid ett enklare sätt att göra det. När man tittar direktpå enkelt sätt, särskilt under långa perioder, du kommer inte att se det.Inte heller kommer Iles.
		-- Rich Hall, "Sniglets"

%
Imbesi lag med Freemans Extension:För att något ska bli ren, något annat måstebli smutsig; men du kan få allt smutsig utan att fånågot ren.
		-- Rich Hall, "Sniglets"

%
Oföränderlighet, tre arbets:(1) Om en presenning kan fladdra, det kommer.(2) Om en liten pojke kan bli smutsig, kommer han.(3) Om en tonåring kan gå ut, kommer han.
		-- Rich Hall, "Sniglets"

%
Opartisk, adj .:Det går inte att uppfatta något löfte av personlig nytta avespousing endera sidan av en kontrovers eller anta någon av tvåmotstridiga åsikter.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
inkorgen, N .:En fångstbassäng för allt du inte vill ta itu med, menär rädda för att kasta bort.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
incitamentsprogram, n .:Systemet med långa och korta belöningar som ett företag användningsområdenatt motivera sitt folk. Fortfarande, trots alla experiment medvinstdelning, aktieoptioner och liknande, det mest effektivaincitamentsprogram hittills verkar vara "Gör ett bra jobb och du får	behåll det."
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kyrkoherdet, n .:Person livligaste intresse för outcumbents.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
index, n .:Alfabetisk lista över ord ingen möjlig intresse där enalfabetisk lista över ämnen med referenser borde vara.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Linda, n .:Perioden av våra liv när, enligt Wordsworth, "Heaven liggerom oss. "Världen börjar ljuga om oss ganska snart efteråt.
		-- Ambrose Bierce

%
Information Center, n .:Ett rum bemannad av professionella dator människor vars jobb det är attberätta varför du inte kan få den information du behöver.
		-- Ambrose Bierce

%
Informationsbearbetning:Vad du kallar databehandling när folk är så äckladdet kommer de inte att låta det att diskuteras i deras närvaro.
		-- Ambrose Bierce

%
Otacksam, n .:En man som biter den hand som föder honom, och sedan klagar övermatsmältningsbesvär.
		-- Ambrose Bierce

%
bläck, n .:En skurkaktig förening tannogallate av järn, gummi arabicum,och vatten, främst för att underlätta infektion avidioti och främja intellektuell brott.
		-- H. L. Mencken

%
förnya, v .:Att irritera folk.
		-- H. L. Mencken

%
osäkerhet, n .:Ta reda på att du har mispronounced för år en av dinafavorit ord.Förverkliga halvvägs genom ett skämt som du säger det tillden person som sa det till dig.
		-- H. L. Mencken

%
intresse, n .:Vilka låntagare betalar, långivare får, aktieägare äger, ochutbrända anställda måste låtsas.
		-- H. L. Mencken

%
Tolk, n .:En som gör det möjligt för två personer av olika språk för attförstå varandra genom att upprepa varje vad det skulle ha varit atttolkens fördel för andra att ha sagt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
berusade, adj .:När du känner sofistikerade utan att kunna uttala det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Iron lag Distribution:Dem som har, blir.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
ISO applikationer:En lösning på jakt efter ett problem!
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Issawi lagar Progress:Jaga av Progress:Det mesta får stadigt värre.Den Path of Progress:En genväg är det längsta avståndet mellan två punkter.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Det är fruktlöst:att bli lachrymose över precipitately avgick laktat vätska.att försöka indoktrinera en avdankad hund medinnovativa manövrar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
"Det är i process":Så insvept i byråkrati att situationen är nästan hopplöst.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
kursiv, adj:Lutar åt höger för att betona nyckelfraser. unikt förVästerländska alfabet; i östra språk, samma fraserofta lutar åt vänster.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Jacquin postulatet om demokratisk regering:Ingen man liv, frihet eller egendom är säkra medanlagstiftaren i sessionen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Jenkinson lag:Det kommer inte att fungera.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Jim Nasium lag:I ett stort omklädningsrum med hundratals skåp, de få människormed hjälp av anläggningen vid någon tidpunkt kommer alla har skåp bredvidvarandra så att alla är trångt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
anställningsintervju, n .:Olidlig process under vilken personaltjänstemänskilja agnarna från vetet - sedan hyra vetet.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
arbetsförmedling, n .:Tala om för din chef vad han kan göra med ditt jobb.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
jogger, n .:En udda slags person med en sak för smärta.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Johnny Carson: s definition:Den minsta tidsintervall som människan känner till är den som skeri Manhattan mellan trafiksignalen bli grönt ochtaxichauffören bakom du blåser hans horn.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Johnsons första lag:När någon mekanisk inrättning misslyckas, kommer den att göra så vidmest obekväma möjliga tid.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Johnsons lag:System liknar de organisationer som skapar dem.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Jones första lag:Den som ger ett betydande bidrag till alla områden försträva, och stannar i detta område tillräckligt länge, blir enobstruktion till dess framsteg - i direkt proportion till denbetydelsen av deras originella bidrag.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Jones Motto:Vänner kommer och går, men fiender ackumuleras.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Jones andra lag:Mannen som ler när saker går fel har tänkt på någonatt skylla det på.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Juall lag om Nice Guys:Trevliga killar inte alltid avsluta sista, ibland inte avsluta.Ibland inte ens får en chans att börja!
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Rättvisa, n .:Ett beslut till din fördel.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Kafkas lag:I kampen mellan dig och världen, tillbaka världen.
		-- Franz Kafka, "RS's 1974 Expectation of Days"

%
Karlson teorem Snack matpaket:För alla P, där P är ett paket med snacks, P är en portionspaket av snacks.Gibson katten Corrolary:För alla L, där L är ett paket med lunch kött, L är Gibson paketlunch kött.
		-- Franz Kafka, "RS's 1974 Expectation of Days"

%
Katz 'lag:Män och nationer kommer att agera rationellt näralla andra möjligheter är uttömda.Historien lär oss att män och nationer beter klokt när de haruttömt alla andra alternativ.
		-- Abba Eban

%
Kaufman första lag Party fysik:Befolkningstätheten är omvänt proportionelltill kvadraten på avståndet från fatet.
		-- Abba Eban

%
Kaufman lag:En policy är en restriktiv dokument för att förhindra en upprepningav en enda incident, där den händelsen aldrig nämns.
		-- Abba Eban

%
Tänk alltid de fyra konstanta lagar Frisbee:(1) Den starkaste kraften i världen är som en skivaansträngande att landa i en bil, precis utom räckhåll (dettakraft är tekniskt kallas "bil suger").(2) föregå aldrig någon manöver av en kommentar mer förutsägandeän "Titta på det här!"(3) Sannolikheten för en frisbee slå något är direktproportionell mot kostnaden för att slå det. Till exempel kan enFrisbee kommer alltid att gå direkt mot en polis elleren gammal dam i stället för beat upp Chevy.(4) Det bästa kast händer när ingen ser; närsöt flicka som du har försökt att imponera tittar, denFrisbee kommer alltid studsa ut din hand eller slå digi huvudet och slå dig dum.
		-- Abba Eban

%
Kennedys Market Sats:Med tanke på tillräckligt insiderinformation och obegränsad kredit,du har att gå sönder.
		-- Abba Eban

%
Kents heuristisk:Leta efter det första där du skulle helst vilja hitta det.
		-- Abba Eban

%
kern, v .:1. För att packa typ tillsammans så tätt som kärnorna på ett öraav majs. 2. I delar av Brooklyn och Queens, NY, en liten,metallföremål som en del av det monetära systemet.
		-- Abba Eban

%
kärna, n .:En del av ett operativsystem som bevarar den medeltidatraditioner trolldom och svart magi.
		-- Abba Eban

%
Kettering Observations:Logic är ett organiserat sätt att gå fel med tillförsikt.
		-- Abba Eban

%
Kime lag för belöning av Ödmjukhet:Vända andra kinden endast ger två blåmärken kinder.
		-- Abba Eban

%
Kin, n .:En åkomma av blodet.
		-- Abba Eban

%
Kington lag för perforering:Om en rak linje av hål görs i en bit papper, såsomsom ett ark av frimärken eller en check, blir den starkaste den linjendelen av pappret.
		-- Abba Eban

%
Kinkler första lag:Ansvaret överstiger alltid myndigheten.Kinkler andra lag:Alla de enkla problem har lösts.
		-- Abba Eban

%
Kliban första lag Mat:äter aldrig något större än ditt huvud.
		-- Abba Eban

%
Kludge, n .:En omaka samling av dåligt matchande delar, som bildar endistressing helhet.
		-- Jackson Granholm, "Datamation"

%
Knebel lag:Det är nu bevisat bortom allt tvivel att rökning är en av de ledandeorsakerna till statistik.
		-- Jackson Granholm, "Datamation"

%
kunskap, n .:Saker du tror.
		-- Jackson Granholm, "Datamation"

%
Kramer lag:Du kan aldrig tala om vilken väg tåget gick genom att titta på spåren.
		-- Jackson Granholm, "Datamation"

%
Krogt, n. (Kemisk beteckning: Kr):Den metalliska silverbeläggning finns på snabbmats spelkort.
		-- Rich Hall, "Sniglets"

%
Labor, n .:En av de processer genom vilka A förvärvar fastighet för B.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Lackland s lagar:(1) aldrig vara först.(2) aldrig vara sist.(3) frivillig aldrig för någonting
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Lactomangulation, n .:Manhandling den "öppna här" pip på en mjölkkartong så illaatt man måste ta till användning av "olaglig" sida.
		-- Rich Hall, "Sniglets"

%
Langsam s lagar:(1) Allt beror på.(2) Ingenting är alltid.(3) Allt är ibland.
		-- Rich Hall, "Sniglets"

%
Larkinson lag:Alla lagar är i grunden falskt.
		-- Rich Hall, "Sniglets"

%
laser, n .:Misslyckades död ray.
		-- Rich Hall, "Sniglets"

%
Lauras lag:Inget barn kastar upp i badrummet.
		-- Rich Hall, "Sniglets"

%
Lagen om kommunikation:Det oundvikliga resultatet av förbättrade och förstorade kommunikationmellan olika nivåer i en hierarki är en kraftigt ökadområde missförstånd.
		-- Rich Hall, "Sniglets"

%
Lagen om Kontinuitet:Experiment bör vara reproducerbar. De bör alla misslyckas på samma sätt.
		-- Rich Hall, "Sniglets"

%
Lagen om förhalning:Förhalning undviker ledan; man aldrig haren känsla av att det inte finns något viktigt att göra.
		-- Rich Hall, "Sniglets"

%
Lagen om Selektiv Gravity:Ett objekt kommer att falla så att göra mest skada.Jenning s Korollarium:Chansen att brödet som faller med den smörade sidanner är direkt proportionell mot kostnaden för mattan.Lagen om perversa naturen:Du kan inte bestämma i förväg vilken sida av bröd smör.
		-- Rich Hall, "Sniglets"

%
Djungelns lag:Den som tvekar är lunch.
		-- Rich Hall, "Sniglets"

%
Laws of Computer Programming:(1) ett visst program, när du kör, är föråldrad.(2) ett visst program kostar mer och tar längre tid.(3) Om ett program är användbar, måste den bytas ut.(4) Om ett program är värdelös, kommer det måste dokumenteras.(5) ett visst program kommer att expandera för att fylla alla tillgängliga minnet.(6) Värdet av ett program är proportionell mot vikten av sin produktion.(7) Program komplexitet växer tills det överskrider kapaciteten hosprogrammeraren som måste behålla den.
		-- Rich Hall, "Sniglets"

%
Lagar Serendipity:(1) För att upptäcka något, måste du vara ute efter något.(2) Om du vill göra en förbättrad produkt, måste du redanatt vara engagerade i en sämre en.
		-- Rich Hall, "Sniglets"

%
stämning, n .:En maskin som du går in som en gris och komma ut som en korv.
		-- Ambrose Bierce

%
Advokat härskar:När lagen är emot dig, hävdar fakta.När fakta är emot dig, hävdar lagen.När båda är emot dig, kallar andra advokat namn.
		-- Ambrose Bierce

%
Lazlo kinesiska Relativity Axiom:Oavsett hur stor din triumfer eller hur tragiskt dina nederlag -cirka en miljard kineser kan inte bry sig mindre.
		-- Ambrose Bierce

%
inlärningskurva, n .:En häpnadsväckande ny teori, upptäcktes av managementkonsulterpå 1970-talet, hävdar att ju mer du gör något somsnabbare du kan göra det.
		-- Ambrose Bierce

%
Lee lag:Mamma sa att det skulle finnas dagar som denna,men hon har aldrig sagt att det skulle vara så många!
		-- Ambrose Bierce

%
Leibowitz härskar:När hamrar på en spik, kommer du aldrig träffa dinfinger om du håller hammaren med båda händerna.
		-- Ambrose Bierce

%
Lemma: Alla hästar har samma färg.Bevis (genom induktion):Fall n = 1: I en uppsättning med endast en häst, är det uppenbart att allahästar i den uppsättningen har samma färg.Fall n = k: Anta att du har en uppsättning av k + 1 hästar. Dra en av dessahästar av den inställda, så att du har k hästar. Antag att allaav dessa hästar har samma färg. Nu sätter tillbaka hästen som dutog ut, och dra ut en annan. Antag att alla de khästar nu i uppsättningen har samma färg. Då uppsättningen k + 1 hästarär alla samma färg. Vi har k sant => k + 1 true; därför allahästar har samma färg.Sats: Alla hästar har ett oändligt antal ben.Bevis (genom hot):Alla håller med om att alla hästar har ett jämnt antal ben. Detär också väl känt att hästar har framben framför och två ben itillbaka. 4 + 2 = 6 ben, som visserligen är ett udda antal ben för enhäst att ha! Nu är det enda nummer som är både jämna och udda äroändlighet; därför alla hästar har ett oändligt antal ben.Emellertid antar att det finns en häst någonstans som inte har enoändligt antal ben. Tja, skulle det vara en häst av en annanfärg; och av Lemma, existerar det inte.
		-- Ambrose Bierce

%
hävstångseffekt, n .:Även om någon inte bry sig om vad världen tyckerom dem, de alltid hoppas att deras mor inte ta reda på.
		-- Ambrose Bierce

%
Lewis lag Travel:Den första delen av bagage ut ur rännan tillhör inte någon,någonsin.
		-- Ambrose Bierce

%
Liar, n .:En advokat med en kringflackande provision.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Lögnare:en som berättar en obehaglig sanning.
		-- Oliver Herford

%
Lie, n .:En mycket dålig ersättning för sanningen, men den endaupptäckts hittills.
		-- Oliver Herford

%
Lieberman lag:Alla ligger, men det spelar ingen roll eftersom ingen lyssnar.
		-- Oliver Herford

%
liv, n .:En infall av flera miljarder celler att vara er för ett tag.
		-- Oliver Herford

%
liv, n .:Lär dig mer om människor den hårda vägen - genom att vara en.
		-- Oliver Herford

%
liv, n .:Det korta mellanspel mellan intighet och evighet.
		-- Oliver Herford

%
fyr, N .:En hög byggnad på stranden där regeringenupprätthåller en lampa och vän av en politiker.
		-- Oliver Herford

%
tycka om:När lever samtidigt är en underbar tillfällighet.
		-- Oliver Herford

%
Linus lag:Det finns ingen tyngre börda än en stor potential.
		-- Oliver Herford

%
Lisp, v .:Om du vill ringa en spade en thpade.
		-- Oliver Herford

%
Lockwood långskott:Chansen att bli uppäten av ett lejon på Main Streetär inte en på miljonen, men en gång skulle vara tillräckligt.
		-- Oliver Herford

%
älskar, n .:Kärleksband i en knut i änden av repet.
		-- Oliver Herford

%
älskar, n .:När det växer, behöver du inte har något emot vattna den med några tårar.
		-- Oliver Herford

%
älskar, n .:När du inte vill att någon alltför nära - att du är mycket känsligtill njutning.
		-- Oliver Herford

%
älskar, n .:När du tänker på någon på dagar som börjar med en morgon.
		-- Oliver Herford

%
älskar, n .:När om han uppmanas att välja mellan din älskareoch lycka, skulle du hoppa lycka i ett pulsslag.
		-- Oliver Herford

%
kärlek, v .:Jag ska låta dig leka med mitt liv om du ska låta mig spela med er.
		-- Oliver Herford

%
Lowery lag:Om det fastnar - tvinga den. Om den går sönder, det behövs ersätter ändå.
		-- Oliver Herford

%
Lubarsky lag av Cybernetic Entomology:Det finns alltid en mer bugg.
		-- Oliver Herford

%
Dårhus, n .:Den plats där optimism mest krusidullar.
		-- Oliver Herford

%
Maskinoberoende, adj .:Inte köras på någon befintlig maskin.
		-- Oliver Herford

%
Mad, adj .:Påverkas med en hög grad av intellektuell självständighet ...
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Madisons Förfrågan:Om du måste resa på Titanic, varför inte gå första klass?
		-- Ambrose Bierce, "The Devil's Dictionary"

%
MAFIA, n:[Förkortning för mekaniserade applikationer tvångs InsuranceRedovisning.] Ett omfattande nätverk med många on-line och off-shoredelsystem som körs under OS, DOS och IOS. MAFIA dokumentation ärganska knapphändiga, och maffian försäljningskontor uppvisar att testyovilja att bona fide undersökningar som är kännetecknande för så många DPoperationer. Från den lilla som sipprat ut, förefaller det som omMAFIA verkar under en icke-standardprotokoll, Omerta, en tystlåtenvariant av SNA, där utökade handslag utför också kompliceradesäkerhetsfunktioner. De kända timesharing aspekterna av MAFIA pekar på enmer än vanligt enväldiga operativsystem. Skärmen bära enimperativ, nonrefusable viktning (de flesta menyer erbjuder enkla JA / JAalternativ, försumliga till YES) som utesluter likgiltighet eller försening.Unikt är all redigering i MAFIA utförs centralt, med hjälp av enkraftfull rubout funktionen kan radera filer, filors, filees, ochhela nodala aggravations.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Magary princip:När det finns en folkstorm för att minska död ved och fett från allastatliga byråkratin, är det död ved och fett som görstyckning och offentliga tjänster skärs.
		-- Stan Kelly-Bootle, "The Devil's DP Dictionary"

%
Magnet, n .:Något som påverkas av magnetism.Magnetism, n .:Något som verkar på en magnet.De två definition omedelbart föregående kondenseras från verk avettusen framstående forskare, som har belysta föremål meden stor vit ljus, till outsägliga utvecklingen av mänsklig kunskap.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Magnocartic, adj .:Alla bil som, när det lämnas obevakat, lockar kundvagnar.
		-- Sniglets, "Rich Hall & Friends"

%
Skata, n .:En fågel vars theivish disposition föreslog någon att detkan läras att prata.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Maier lag:Om fakta inte överensstämmer med teorin, måste de tas om hand.korollarier:(1) Ju större teorin, desto bättre.(2) Experimentet kan betraktas som en framgång om inte mer än50% av de observerade mätningarna måste kasseras tillerhålla en korrespondens med teorin.
		-- N. R. Maier, "American Psychologist", March 1960

%
Huvud lag:För varje handling finns en likvärdig och motsatt regeringsprogrammet.
		-- N. R. Maier, "American Psychologist", March 1960

%
Ansvarig motto:Om vi ​​inte kan fixa det, är det inte bröt.
		-- N. R. Maier, "American Psychologist", March 1960

%
Major premiss:Sextio män kan göra sextio gånger så mycket arbete som en människa.Mindre premiss:En man kan gräva en Stolphål i sextio sekunder.Slutsats:Sextio män kan gräva en Stolphål i en sekund.Sekundär Slutsats:Inser du hur många hål det skulle vara om folkskulle bara ta sig tid att ta smuts borta från dem?
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Majoriteten, n .:Att kvalitet som skiljer ett brott från en lag.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Man, n .:En medlem av ogenomtänkta eller försumbar kön. Hanen avmänskligheten är allmänt känt att den kvinnliga som Mere Man. släktethar två varianter: bra leverantörer och dåliga leverantörer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Malek lag:Någon enkel idé kommer att formuleras i det mest komplicerade sätt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
felbehandling, n .:Anledningen kirurger bär masker.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
ledning, n .:Konsten att få andra människor att göra allt arbete.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
manodepressiv, adj .:Lätt glum, lätt glöd.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Manlys Maxim:Logik är en systematisk metod för att komma till fel slutsatser	med självförtroende.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
manual, n .:En enhet av dokumentation. Det finns alltid tre eller mer på en vissobjekt. En är på hyllan; någon har de andra. Informationendu behöver finns i de andra.
		-- Ray Simard

%
Marks Dental ordförande Discovery:Tandläkare är oförmögna att ställa frågor som kräver enenkelt ja eller nej.
		-- Ray Simard

%
äktenskap, n .:En gammal, etablerad institution, som ingås mellan två personer djupti kärlek och önskar att göra en engagemang för varandra uttryckaden kärleken. Kort sagt, engagemang för en institution.
		-- Ray Simard

%
äktenskap, n .:Konvertibla obligationer.
		-- Ray Simard

%
Förbindelse, n .:Den onda aye.
		-- Ray Simard

%
Marxistiska lagen om fördelning av välståndet:Brist kommer att delas lika mellan bönderna.
		-- Ray Simard

%
Maryann lag:Du kan alltid hitta det du inte är ute efter.
		-- Ray Simard

%
Maslows Maxim:Om det enda verktyg man har är en hammare, behandlar dig allt somen spik.
		-- Ray Simard

%
Mason första lag Synergism:En dag du vill sälja din själ för något, själar är ett överflöd.
		-- Ray Simard

%
matematiker, n .:Någon som tror imaginära saker att visa sig innan _ i talet.
		-- Ray Simard

%
Matz lag:En slutsats är den plats där du tröttnade att tänka.
		-- Ray Simard

%
Maj lag:Kvaliteten på korrelationen är inversly proportionell mot densitetenav kontroll. (Ju färre datapunkter, desto jämnare kurvorna.)
		-- Ray Simard

%
McEwan härskar av relativa betydelse:När du reser med en besättning av elefanter, inte vara den första attligga ner och vila.
		-- Ray Simard

%
McGowan Madison Avenue Axiom:Om ett objekt marknadsförs som "under $ 50", kan du satsa det är inte $ 19.95.
		-- Ray Simard

%
Meade Maxim:Alltid komma ihåg att du är helt unik, precis som alla andra.
		-- Ray Simard

%
Meader lag:Vad som än händer dig, det kommer tidigarehar hänt med alla du känner, bara mer så.
		-- Ray Simard

%
möte, n .:En sammansättning av människor som kommer samman för att bestämma vilken person elleravdelning som inte är representerad i rummet måste lösa ett problem.
		-- Ray Simard

%
möten, n .:En plats där minuter hålls och timmar förlorade.
		-- Ray Simard

%
memo, n .:Ett interoffice kommunikation alltför ofta skrivit mer till förmånav den person som skickar det än den person som tar emot det.
		-- Ray Simard

%
Mencken och Nathans femtonde lag den genomsnittlige amerikanen:Den värsta skådespelerska i bolaget är alltid chefens fru.
		-- Ray Simard

%
Mencken och Nathan nionde lag den genomsnittlige amerikanen:Kvaliteten på en champagne bedöms av mängden bullerkork gör när den är poppade.
		-- Ray Simard

%
Mencken och Nathans andra lag den genomsnittlige amerikanen:Alla postmästare i småstäder läst alla vykort.
		-- Ray Simard

%
Mencken och Nathans sextonde lag den genomsnittlige amerikanen:Mjölka en ko är en operation som kräver en speciell talang somär besatt endast lantisarna, och ingen person är född i en storstad kannågonsin hoppas att få det.
		-- Ray Simard

%
Meny, n .:En lista över rätter som restaurangen bara har slut på.
		-- Ray Simard

%
Meskimen lag:Det finns aldrig tid att göra det rätt, men det finns alltid tid attgöra det över.
		-- Ray Simard

%
meterologist, n .:Den som tvivlar på etablerat faktum att det ärskyldig att regna om du glömmer ditt paraply.
		-- Ray Simard

%
Mikro Credo:Aldrig lita på en dator större än du kan lyfta.
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
micro:Tänkare leksaker.
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
Miksch lag:Om en sträng har en ände, då har det en annan ände.
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
Miller slogan:Förlora några, förlorar några.
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
millihelen, n .:Mängden av skönhet som krävs för att lansera ett skepp.
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
minidator:En dator som kan ges på budgeten för ett medelnivå manager.
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
MIPS:Menings indikatorn för processorhastighet
		-- Mrs. Byrne's Dictionary of Unusual, Obscure, and

%
Olycka, n .:Den typ av förmögenhet som aldrig missar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
MIT:Georgia Tech i norr
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Mitchell lag av kommittéer:Alla enkla problem kan göras olöslig om tillräckligt många mötenför att diskutera det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
mittsquinter, adj .:En basebollspelare som ser in i hans handske efter att ha missat bollen, somom, på något sätt, orsaken till felet ligger där.
		-- "Sniglets", Rich Hall & Friends

%
Mix lag:Det finns inget mer permanent än en tillfällig byggnad.Det finns inget mer permanent än en tillfällig skatt.
		-- "Sniglets", Rich Hall & Friends

%
blandade känslor:Titta på en busslast med advokater störta från en klippa.Med fem tomma platser.
		-- "Sniglets", Rich Hall & Friends

%
blandade känslor:Titta på din mamma-in-law tillbaka från en klippa ...i ditt nya Mercedes.
		-- "Sniglets", Rich Hall & Friends

%
modem, adj .:Up-to-date, nymodig, som i "Grundligt Modem Millie." Enolycklig biprodukt av kerning.[Det är sic!]
		-- "Sniglets", Rich Hall & Friends

%
blygsamhet, n .:Vara bekväm att andra kommer att upptäcka din storhet.
		-- "Sniglets", Rich Hall & Friends

%
Anspråkslöshet:Den milda konsten att förbättra din charm genom att låtsas att inte varamedvetna om det.
		-- Oliver Herford

%
Molekyl, n .:Den ultimata, odelbar enhet materia. Men är inte detsammafrån blodkropp, även den ultimata, odelbar enhet materia, genom ennärmare likhet med atomen, också det ultimata, odelbar enhetmateria ... Jon skiljer sig från molekylen, den blodkropp ochatomen i att det är en jon ...
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Mollison byråkrati Hypotes:Om en idé kan överleva en byråkratisk översyn och genomförasdet var inte värt att göra.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
fart, n .:Vad du ge en person när de går bort.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Moon, n .:1. En himlakropp vars fas är mycket viktigt för hackare. SeMånfas. 2. Dave månen (MOON @ MC).
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Moores konstant:Alla syftar till att göra något, och allagör något, men ingen gör vad han syftar till att göra.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
mophobia, n .:Rädsla för att bli muntligen missbrukas av en Mississippian.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Morton lag:Om råttor experimenterat på, kommer de att utveckla cancer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Mosher lag för programvaruteknik:Oroa dig inte om det inte fungerar rätt. Om allt gjorde, skulle duvara utan jobb.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Mr Coles Axiom:Summan av intelligens på planeten är en konstant; debefolkningen växer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
mamma, n .:En egyptier som var ont om tid.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Murphys lag för forskning:Nog forskning tenderar att stödja din teori.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Murphys lagar:(1) Om något kan gå fel, kommer det.(2) Ingenting är så lätt som det ser ut.(3) Allt tar längre tid än du tror att det kommer.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Murrays Regel:Varje land med "demokratiska" i titeln är inte.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Mustgo, n .:Någon del av mat som har suttit i kylskåpet sålänge har det blivit ett forskningsprojekt.
		-- Sniglets, "Rich Hall & Friends"

%
Min far lärde mig tre saker:(1) Blanda aldrig whisky med något annat än vatten.(2) Försök aldrig att dra till en hålstege.(3) diskutera aldrig affärer med någon som vägrar att ge sitt namn.
		-- Sniglets, "Rich Hall & Friends"

%
Nachman härskar:När det gäller utländsk mat, desto mindre autentiska desto bättre.
		-- Gerald Nachman

%
narcolepulacyi, n .:Den smittsamma verkan gäspningar, vilket alla i sikteockså gäspning.
		-- "Sniglets", Rich Hall & Friends

%
nerd pack, n .:Plastficka bärs i bröstfickan för att hålla pennor från nedsmutsningkläder. Nerd position inom teknik hierarkin kan mätasgenom antalet pennor, fett pennor och linjaler bristling i sin förpackning.
		-- "Sniglets", Rich Hall & Friends

%
neutron bomb, n .:En sprängladdning av begränsat militärt värde eftersom, somdet bara förstör människor utan att förstöra egendom, detmåste användas tillsammans med bomber som förstör egendom.
		-- "Sniglets", Rich Hall & Friends

%
nytt, adj .:Annan färg än tidigare modell.
		-- "Sniglets", Rich Hall & Friends

%
Newlan s Truism:En "acceptabel" nivå av arbetslöshet innebär attregering ekonom som det är acceptabelt fortfarande har ett jobb.
		-- "Sniglets", Rich Hall & Friends

%
Newman Discovery:Din bästa drömmar kan inte gå i uppfyllelse; lyckligtvis, inte heller kommerdin värsta drömmar.
		-- "Sniglets", Rich Hall & Friends

%
Newtons gravitationslag:Vad går upp måste komma ner. Men förvänta dig inte att komma ner därdu kan hitta den. Murphys lag gäller Newtons.
		-- "Sniglets", Rich Hall & Friends

%
Newtons föga kända sjunde lag:En fågel i handen är säkrare än en overhead.
		-- "Sniglets", Rich Hall & Friends

%
Nick den grekiska lag of Life:Allt som allt är livet 9-5 mot.
		-- "Sniglets", Rich Hall & Friends

%
Ninety-Ninety Rule of Project scheman:Den första nittio procent av uppgiften tar nittio procent avtiden, och den sista tio procent tar den andra nittio procent.
		-- "Sniglets", Rich Hall & Friends

%
enkel:Ett beslut som, sedd genom retrospectoscope,är "uppenbart" till dem som inte gör det från början.
		-- "Sniglets", Rich Hall & Friends

%
inget underhåll:Omöjligt att fastställa.
		-- "Sniglets", Rich Hall & Friends

%
nolo contendere:En juridisk term som betyder: "Det var inte jag, domare, och jag kommer aldrig att göra	det igen."
		-- "Sniglets", Rich Hall & Friends

%
nominell ägg:Nya Yorkerese för dyra.
		-- "Sniglets", Rich Hall & Friends

%
Ensidiga lagar Förväntningarna:Negativa förväntningar ger negativa resultat.Positiva förväntningar ger negativa resultat.
		-- "Sniglets", Rich Hall & Friends

%
Nouvelle cuisine, n .:Franska för "inte tillräckligt med mat".Kontinental frukost, n .:Engelska för "inte tillräckligt med mat".Tapas, n .:Spanska för "inte tillräckligt med mat".Dim Sum, n .:Kinesiska för mer mat än du någonsin sett i hela ditt liv.
		-- "Sniglets", Rich Hall & Friends

%
November, n .:Den elfte tolftedel av en trötthet.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Novinson revolutionära Discovery:När kommer revolutionen, kommer saker och ting att vara annorlunda -inte bättre, bara annorlunda.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Nowlan teori:Den som tvekar är inte bara förlorat, men flera miles frånnästa avfart motorväg.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Nusbaum härskar:Ju mer pretentiös den firma, ju mindreorganisation. (Till exempel Murphy centret förKodifiering av mänskliga och organisatoriska lag, kontrasteIBM, GM, och AT & T.)
		-- Ambrose Bierce, "The Devil's Dictionary"

%
O'Brian lag:Allt sker alltid av fel skäl.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
O'Reilly lag av kök:Renlighet är näst intill omöjligt
		-- Ambrose Bierce, "The Devil's Dictionary"

%
O'Toole s kommentar till Murphys lag:Murphy var en optimist.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Occams suddgummi:Den filosofiska principen att även den enklasteLösningen är skyldig att ha något fel med det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Office Automation:Användningen av datorer för att förbättra effektiviteten på kontoretgenom att ta bort någon du skulle vilja prata med över kaffe.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Officiella projektfaser:(1) okritiskt accepterande(2) Wild Entusiasm(3) nedslagen Disillusionment(4) total förvirring(5) Sök efter den Guilty(6) bestraffning av oskyldiga(7) Främjande av icke-deltagare
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ogden lag:Ju tidigare du halkar efter, desto mer tid du har att komma ikapp.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Gammalt japanskt ordspråk:Det finns två typer av dårar - de som aldrig klättra Mt. Fuji,och de som klättrar den två gånger.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Gammal tidmätare, n .:En som minns när välgörenhet var en dygd och inte en organisation.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Oliver lag:Erfarenhet är något du inte får förrän strax efter att du behöver det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Olmstead lag:När allt är sagt och gjort, är en fan av mycket mer sagt än gjort.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
omnibiblious, adj .:Likgiltig för typ av dryck. Ex: "Åh, du kan få mig något.Jag omnibiblious. "
		-- Ambrose Bierce, "The Devil's Dictionary"

%
På förmåga:En dvärg är liten, även om han står på en bergstopp,en koloss håller sin höjd, även om han står i en brunn.
		-- Lucius Annaeus Seneca, 4BC - 65AD

%
När det gäller C-program indrag:"I min Egotistical yttrande, bör de flesta människors C-program varaindragen sex fot nedåt och täckt med smuts. "
		-- Blair P. Houghton

%
On-line, adj .:Tanken att en människa ska alltid vara tillgängliga för en dator.
		-- Blair P. Houghton

%
En gång, adv .:	Tillräckligt.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
One Page Princip:En specifikation som inte får plats på en sida av 8,5x11 tumpapper kan inte förstås.
		-- Mark Ardis

%
"En storlek passar alla":Passar inte någon.
		-- Mark Ardis

%
One Shot Fallstudie, n .:Den vetenskapliga ekvivalent av klöver fyra blad, från vilken det ärslutsatsen alla klöver har fyra blad och ibland grönt.
		-- Mark Ardis

%
Optimism, n .:Tron att allt är vacker, inklusive vad som är fult, bra,dålig, och allt rätt som är fel. Den hålls med störstuthållighet av dem vana vid att falla i motgångar, och de flestaacceptabelt framförts med flin som aporna ett leende. Som en blindtro, är den oåtkomlig för ljuset av motbevis - en intellektuelloordning, vilket ger ingen behandling men död. Det är ärftlig, meninte smittsam.
		-- Mark Ardis

%
optimist, n .:En förespråkare av den uppfattningen att svart är vitt.En pessimist bad Gud om hjälp."Ah, du vill mig att återställa hopp och glädje", säger Gud."Nej", svarade framställaren, "Jag önskar dig att skapa något somskulle motivera dem. ""Världen är alla skapade," sade Gud, "men du har förbisettnågot - dödligheten av optimisten ".
		-- Ambrose Bierce, "The Devil's Dictionary"

%
optimist, n:En säckpipor med en personsökare.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Oregano, n .:Den antika italienska konsten pizza vikning.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Osborn lag:Variabler inte; konstanter är inte.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ozman s lagar:(1) Om någon säger att han kommer att göra något "utan att misslyckas", han kommer inte.(2) Ju fler människor talar i telefon, desto mindre pengar de gör.(3) Människor som går till konferenser är de som inte borde.(4) Pizza brinner alltid gommen.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
smärta, n .:En sak, åtminstone det visar sig att du lever!
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Målning, n .:Konsten att skydda plana ytor från väder ochutsätta dem för kritikern.
		-- Ambrose Bierce

%
Pandoras Regel:Öppna aldrig en låda du inte stänga.
		-- Ambrose Bierce

%
Paprika Åtgärd:2 streck == 1 smidgen2 smidgens == en nypa3 krm == en Soupcon2 soupcons == 2 mycket paprika
		-- Ambrose Bierce

%
paranoia, n .:En hälsosam förståelse för hur universum fungerar.
		-- Ambrose Bierce

%
Pardo första postulat:Något bra i livet är antingen olagligt, omoraliskt, eller gödning.Arnolds Addendum:Allt annat orsakar cancer hos råttor.
		-- Ambrose Bierce

%
Parkinsons femte lag:Om det finns ett sätt att fördröja i viktiga beslut, det godabyråkrati, offentlig eller privat, kommer att finna det.
		-- Ambrose Bierce

%
Parkinsons fjärde lag:Antalet personer i någon arbetsgrupp tenderar att ökaoavsett hur mycket arbete som skall utföras.
		-- Ambrose Bierce

%
parti, N .:En samling där du möter människor som drickerså mycket du kan inte ens komma ihåg deras namn.
		-- Ambrose Bierce

%
Pascal Användare:Pascal-systemet kommer att ersättas nästa tisdag med Cobol.Ändra dina program i enlighet med detta.
		-- Ambrose Bierce

%
Pascal Användare:För att visa respekt för 313th årsdag (i morgon) idöd Blaise Pascal, kommer dina program att köras på halvfart.
		-- Ambrose Bierce

%
Pascal:Ett programmeringsspråk uppkallad efter en man som skulle vändai sin grav om han visste om det.
		-- Datamation, January 15, 1984

%
Lösenord:
		-- Datamation, January 15, 1984

%
Patageometry, n .:Studien av de matematiska egenskaper som är invariantenligt hjärntransplantat.
		-- Datamation, January 15, 1984

%
patent:En metod för att sprida uppfinningar så att andra kan kopiera dem.
		-- Datamation, January 15, 1984

%
Paul lag:I Amerika, det är inte hur mycket en artikelkostnader, det är hur mycket du sparar.
		-- Datamation, January 15, 1984

%
Paul lag:Du kan inte falla från golvet.
		-- Datamation, January 15, 1984

%
lön:Den veckovisa $ 5,27 som återstår efter avdrag för federalakällskatt, statliga källskatt, stad källskatt, FICA,Medicin / tandvård, långvarig arbetsoförmåga, arbetslöshetsförsäkring,Christmas Club, och löne sparplan bidrag.
		-- Datamation, January 15, 1984

%
Fred, n .:I internationella frågor, en period av fusk mellan tvåperioder av strider.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Pecor hälsa-Food Princip:Ät aldrig kålrot på någon dag i veckan som har ett "y" i det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Pedaeration, n .:Den perfekta kroppsvärme uppnås genom att ha ett ben underark och en hängande över kanten på sängen.
		-- Rich Hall, "Sniglets"

%
pediddel:En bil med endast en arbetsdag framlykta.
		-- "Sniglets", Rich Hall & Friends

%
Klienter lag:Lösningen på ett problem förändrar problemets natur.
		-- "Sniglets", Rich Hall & Friends

%
Penguin Trivia # 46:Djur som inte pingviner kan bara önskar att de var.
		-- Chicago Reader 10/15/82

%
pension:En federalt försäkrade kedjebrev.
		-- Chicago Reader 10/15/82

%
Människors Action Regler:(1) En del människor som kan, bör inte.(2) Vissa personer som bör inte.(3) En del människor som inte borde, kommer.(4) En del människor som inte kan, kommer att försöka, oavsett.(5) Vissa människor som borde inte, men försök, kommer då att skylla på andra.
		-- Chicago Reader 10/15/82

%
perfekt gäst:En som gör sin värd känna sig hemma.
		-- Chicago Reader 10/15/82

%
Prestanda:Ett uttalande av den hastighet med vilken ett datorsystem fungerar. Ellersnarare kan fungera under vissa omständigheter. Eller sadesatt arbeta under i Jersey ungefär en månad sedan.
		-- Chicago Reader 10/15/82

%
pessimist:En man som tillbringar all sin tid på att oroa hur han kan hållawolf från dörren.optimist:En man som vägrar att se vargen tills han griper sätebyxorna.opportunistisk:En man som bjuder vargen in och visas nästa dag i en päls.
		-- Chicago Reader 10/15/82

%
Peter lag substitutions:Titta efter mullvadshögar, ochberg kommer att se efter sig själva.Peter Principen om framgång:Få upp en gång mer än du nedslagen.
		-- Chicago Reader 10/15/82

%
Peterson förmaning:När du tror att du kommer ner för tredje gången -bara ihåg att du kan ha räknat fel.
		-- Chicago Reader 10/15/82

%
Peterson regler:(1) Lastbilar som välter på motorvägar är fyllda med något klibbig.(2) Ingen söt baby i en vagn är alltid en flicka när kallas en.(3) Saker som fästing är inte alltid klockor.(4) Självmord fungerar bara när du bluffar.
		-- Chicago Reader 10/15/82

%
petribar:Alla solblekt förhistoriska godis som har suttit ifönstret i en varuautomat för lång.
		-- Rich Hall, "Sniglets"

%
Faser av ett projekt:(1) Exultation.(2) disenchantment.(3) Förvirring.(4) Sök efter de skyldiga.(5) straff för Innocent.(6) Godkänd på oengagerade.
		-- Rich Hall, "Sniglets"

%
filosofi:Förmågan att bära med lugn olyckor av våra vänner.
		-- Rich Hall, "Sniglets"

%
filosofi:Obegripliga svar på olösliga problem.
		-- Rich Hall, "Sniglets"

%
phosflink:Att bläddra en glödlampa på och av när den har brunnit ut (som om något, attkommer att föra den tillbaka till livet).
		-- "Sniglets", Rich Hall & Friends

%
Pickle lag:Om kongressen måste göra en smärtsam sak,saken måste göras i ett udda-antal år.
		-- "Sniglets", Rich Hall & Friends

%
pixel, n .:En busig, magisk anda i samband med skärmar.Datorindustrin har ofta lånat från mytologin:Bevittna sprites i datorgrafik, demonerna inom artificiellintelligens, och trollen på marknadsavdelningen.
		-- "Sniglets", Rich Hall & Friends

%
Notera att:
		-- "Sniglets", Rich Hall & Friends

%
Pohl lag:Ingenting är så bra att någon, någonstans, kommer inte hata det.
		-- "Sniglets", Rich Hall & Friends

%
förgiftat kaffe, n .:Grunder för skilsmässa.
		-- "Sniglets", Rich Hall & Friends

%
politik, n .:En strid intressemaskerats som en tävling av principer.Genomförandet av offentliga angelägenheter för privat fördel.
		-- Ambrose Bierce

%
Pollyanna Educational konstant:Den hyperaktiva barn är aldrig frånvarande.
		-- Ambrose Bierce

%
polygon:Död papegoja.
		-- Ambrose Bierce

%
Poorman härskar:När du drar en plast skräp väska från dess praktiska dispenser paket,du alltid få tag på den slutna änden och försöka dra den öppna.
		-- Ambrose Bierce

%
Bärbar, adj .:Lever omstart.
		-- Ambrose Bierce

%
Positiv, adj .:Misstas på toppen av en röst.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
fattigdom, n .:En olycklig tillstånd som kvarstår så längesom alla saknar något han skulle vilja ha.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ström, n .:Den enda narkotiska regleras av SEC i stället för FDA.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
prärier, n .:Vidsträckta slätter som omfattas av trädlösa skogar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Fördom:En lösdrivare yttrande utan synliga försörjning.
		-- Ambrose Bierce

%
Preudhomme lag av Fönsterputsning:Det är på den andra sidan.
		-- Ambrose Bierce

%
Pris råd:Det är ett spel - spela det att ha kul.
		-- Ambrose Bierce

%
Prioritet:Ett uttalande om vikten av en användare eller ett program. Oftauttryckt som en relativ prioritet, vilket indikerar att användaren intevård när arbetet är slutfört så länge han behandlas mindredåligt än någon annan.
		-- Ambrose Bierce

%
problem dricker, n .:En man som aldrig köper.
		-- Ambrose Bierce

%
programmet, n .:En magisk spell kasta över en dator som gör det möjligt att vända en ingångi felmeddelanden. tr.v. Att engagera sig i ett tidsfördriv som liknar nävenhuvudet mot en vägg, men med färre möjligheter till belöning.
		-- Ambrose Bierce

%
programmet, n .:Varje uppgift som inte kan fyllas i på ett telefonsamtal eller ettdag. När en uppgift definieras som ett program ( "träningsprogram","Försäljningsprogram" eller "marknadsföring programmet"), dess genomförandealltid motiverar att anställa åtminstone ytterligare tre personer.
		-- Ambrose Bierce

%
Programmering Avdelning:Misstag görs medan du väntar.
		-- Ambrose Bierce

%
framsteg, n .:Medeltida man trodde sjukdom orsakades av osynliga demonerinvaderar kroppen och tar i besittning.Den moderna människan vet Sjukdomen orsakas av mikroskopiska bakterieroch virus invaderar kroppen och orsakar det att fungera.
		-- Ambrose Bierce

%
Bevis tekniker # 2: Bevis av Oddity.PROV: För att bevisa att hästar har ett oändligt antal ben.(1) Hästar har ett jämnt antal ben.(2) De har två ben på baksidan och frambenen framför.(3) Detta ger totalt sex ben, vilket säkerligen är ett udda antal    ben för en häst.(4) Men det enda numret som är både udda och jämna är oändligheten.(5) Därför måste hästar ha ett oändligt antal ben.Ämnen är täckas i kommande nummer innehålla bevis efter:skrämselGesticulation (handwaving)"Prova, det fungerar"Förstoppning (jag var bara sitter där och ...)uppenbar påståendeÄndra samtliga 2-talet till _ n s	SamtyckeAvsaknad av ett motexempel, och"Det är självklart"
		-- Ambrose Bierce

%
prototyp, n .:Första steget i livscykeln för en datorprodukt, följt avpre-alfa, alfa, beta, versionen, korrigerad versionen,uppgradera, korrigerad uppgradering, etc. Till skillnad från dess efterföljare, denprototyp förväntas inte att fungera.
		-- Ambrose Bierce

%
Pryor Observations:Hur länge du lever har inget att göramed hur länge du kommer att vara död.
		-- Ambrose Bierce

%
Pudder lag:Allt som börjar väl kommer att sluta illa.(OBS: Det omvända av Pudder lag är inte sant.)
		-- Ambrose Bierce

%
purpitation, n .:Att ta något utanför livsmedelshyllan, bestämmer digvill inte ha det, och sedan lägga den i en annan del.
		-- "Sniglets", Rich Hall & Friends

%
Putt lag:Teknik domineras av två typer av människor:De som förstår vad de inte lyckas.De som lyckas vad de inte förstår.
		-- "Sniglets", Rich Hall & Friends

%
QOTD:"Det är inte förtvivlan ... jag kan stå förtvivlan. Det är hopp."
		-- "Sniglets", Rich Hall & Friends

%
QOTD:"Ett barn av fem kunde förstå detta! Hämta mig ett barn av 5."
		-- "Sniglets", Rich Hall & Friends

%
QOTD:"En universitetsfakultet är 500 egoister med gemensam parkering problem."
		-- "Sniglets", Rich Hall & Friends

%
QOTD:"Luktar du något brännande eller är det mig?"
		-- Joan of Arc

%
QOTD:"Låt inte ditt sinne vandra - det är för lite att släppa ut ensam."
		-- Joan of Arc

%
QOTD:"East är öst ... och låt oss hålla det på det sättet."
		-- Joan of Arc

%
QOTD:"Även Frihetsgudinnan rakar sina gropar."
		-- Joan of Arc

%
QOTD:"Varje morgon jag läsa döds, om mitt namn inte finns där,	Jag går till jobbet."
		-- Joan of Arc

%
QOTD:"Allt jag är idag jag är skyldig till folk, som det är nuför sent att straffa. "
		-- Joan of Arc

%
QOTD:"Han äter som en fågel ... fem gånger sin egen vikt varje dag."
		-- Joan of Arc

%
QOTD:"Han är på samma buss, men han är säker på som fan fick en annanbiljett. "
		-- Joan of Arc

%
QOTD:"Jag inte är trasigt, men jag är dåligt böjd."
		-- Joan of Arc

%
QOTD:"Jag är inte säker på vad det är, men ett" F "skulle bara dignify det."
		-- Joan of Arc

%
QOTD:"Jag tror inte att de skulle kunna sätta honom på ett mentalsjukhus. Påandra sidan, om han redan var i, jag tror inte att de skulle låta honom. "
		-- Joan of Arc

%
QOTD:"Jag kör min bil tyst, för det är självklart."
		-- Joan of Arc

%
QOTD:"Jag har inte kommit tillräckligt långt, och inte kalla mig baby."
		-- Joan of Arc

%
QOTD:"Jag kanske inte kan gå, men jag kör från sittande ställning."
		-- Joan of Arc

%
QOTD:"Jag har aldrig träffat en man som jag inte kunde dricka vacker."
		-- Joan of Arc

%
QOTD:"Jag rör bara bas med verkligheten på ett behov när det behövs!"
		-- Joan of Arc

%
QOTD:"Jag stänkte bakpulver över ett par potatis, men detfungerade inte. "
		-- Joan of Arc

%
QOTD:"Jag trodde att jag såg en enhörning på vägen över, men det var bara enhäst med ett av hornen avbrutna. "
		-- Joan of Arc

%
QOTD:"Jag försökte köpa en get i stället för en trädgårdstraktor, var tvungen att återvändadet dock. Det gick inte att räkna ut ett sätt att ansluta snöslungan. "
		-- Joan of Arc

%
QOTD:"Jag brukade vara en idealist, men jag fick rånad av verkligheten."
		-- Joan of Arc

%
QOTD:"Jag brukade gå förlorad i shuffle, nu jag bara blanda tillsammans med	den försvunna."
		-- Joan of Arc

%
QOTD:"Jag brukade få hög på livet, men på sistone har jag byggt upp ett motstånd."
		-- Joan of Arc

%
QOTD:"Jag brukade gå till UCLA, men sedan min pappa fick ett jobb."
		-- Joan of Arc

%
QOTD:"Jag brukade jogga, men isen höll studsar ut ur mitt glas."
		-- Joan of Arc

%
QOTD:"Jag kommer inte att säga att han är osant, men hans fru har att ringahund för middag. "
		-- Joan of Arc

%
QOTD:"Jag skulle aldrig gifta sig med en kvinna som inte gillar pizza ... Jag kan spelagolf med henne, men jag skulle inte gifta sig med henne! "
		-- Joan of Arc

%
QOTD:"Jag ska ta reson när det kommer ut på CD."
		-- Joan of Arc

%
QOTD:"Jag är bara en pojke som heter" SU "..."
		-- Joan of Arc

%
QOTD:"Jag är inte riktigt för apati, men jag är inte emot det heller ..."
		-- Joan of Arc

%
QOTD:"Jag är på en fisk och skaldjur diet - Jag ser mat och jag äter det."
		-- Joan of Arc

%
QOTD:"Jag har alltid velat arbeta i Förbunds Mint. Och sedan gå vidarestrejk. För att göra mindre pengar. "
		-- Joan of Arc

%
QOTD:"Jag har en sista sak att säga innan jag går, ge mig tillbakaalla mina grejer. "
		-- Joan of Arc

%
QOTD:"Jag har precis lärt om sin sjukdom. Låt oss hoppas att det är ingentingtrivialt. "
		-- Joan of Arc

%
QOTD:"Om han lär sig av sina misstag, ganska snart han vet allt."
		-- Joan of Arc

%
QOTD:"Om jag kunde gå på det sättet, skulle jag inte behöva Köln, nu skulle jag?"
		-- Joan of Arc

%
QOTD:"Om jag vad jag äter, jag är en chocolate chip cookie."
		-- Joan of Arc

%
QOTD:"Om du håller ett öppet sinne folk kommer att kasta en massa skräp i det."
		-- Joan of Arc

%
QOTD:"I köpcentrum i sinnet, är han i leksaksavdelningen."
		-- Joan of Arc

%
QOTD:"Det förefaller mig som antennen inte ta in för mångastationer längre. "
		-- Joan of Arc

%
QOTD:"Det var så kallt i vintras att jag såg en advokat med hanshänderna i egna fickor. "
		-- Joan of Arc

%
QOTD:"Det skulle inte ha varit något, även om det kommer att bli en sak."
		-- Joan of Arc

%
QOTD:"Det är en kall skål med chili, när kärleken inte fungerar."
		-- Joan of Arc

%
QOTD:"Det har varit Måndag hela veckan i dag."
		-- Joan of Arc

%
QOTD:"Det har varit äkta och det har varit kul, men det har inte varit riktigt roligt."
		-- Joan of Arc

%
QOTD:"Det är svårt att säga om han har ett ess i rockärmen eller omess saknas hans däck helt och hållet. "
		-- Joan of Arc

%
QOTD:"Det är en slags hot, du ser. Jag har aldrig varit mycket bra pådem själv, men jag får höra att de kan vara mycket effektivt. "
		-- Joan of Arc

%
QOTD:"Hur mycket kan jag komma undan med och fortfarande komma till himlen?"
		-- Joan of Arc

%
QOTD:"Brist på planering från din sida inte, utgöra en nödsituationfrån min sida. "
		-- Joan of Arc

%
QOTD:"Gillar du ros, kommer vår kärlek vissna och dö."
		-- Joan of Arc

%
QOTD:"Mitt liv är en såpopera, men vem som får filmrättigheterna?"
		-- Joan of Arc

%
QOTD:"Min schampo varar längre än mina relationer."
		-- Joan of Arc

%
QOTD:"Självklart är det mordvapnet. Vem skulle rama in någon med	en falsk?"
		-- Joan of Arc

%
QOTD:"Naturligtvis finns det ingen anledning till det, det är bara vår politik."
		-- Joan of Arc

%
QOTD:"Åh, nej, nej ... Jag är inte vacker. Bara mycket, mycket vacker."
		-- Joan of Arc

%
QOTD:"Våra föräldrar var aldrig vår ålder."
		-- Joan of Arc

%
QOTD:"Övervikt är när du kliver på hundens svans och det dör."
		-- Joan of Arc

%
QOTD:"Säg, du ser ganska atletisk. Vad säger vi sätta ett par tennisskor på dig och kör dig in i väggen? "
		-- Joan of Arc

%
QOTD:"Hon är ungefär lika smart som bete."
		-- Joan of Arc

%
QOTD:"Visst, vände jag ner en drink en gång. Förstod inte frågan."
		-- Joan of Arc

%
QOTD:"Barnet var så ful att de var tvungna att hänga en fläskkotlett runt desshals för att få hunden att leka med den. "
		-- Joan of Arc

%
QOTD:"De äldre gudarna gick till Suggoth och allt jag fick var denna nedlusade T-tröja."
		-- Joan of Arc

%
QOTD:"Det kan inte finnas någon ursäkt för lättja, men jag är säker på att titta."
		-- Joan of Arc

%
QOTD:"Detta är en linje bevis ... om vi börjar tillräckligt långt för att det	vänster."
		-- Joan of Arc

%
QOTD:"Otur? Om jag köpte en pumpa gård, de skulle avbryta Halloween."
		-- Joan of Arc

%
QOTD:"Vad menar du, du hade hunden fast? Precis vad gjorde dutror att han var bruten! "
		-- Joan of Arc

%
QOTD:"Vad jag gillar mest om mig själv är att jag är så förståendeNär jag röra upp saker. "
		-- Joan of Arc

%
QOTD:"Vad kvinnor och psykologer kallar 'släppa din rustning", kallar vi"Blottar halsen."
		-- Joan of Arc

%
QOTD:"När hon halade ass, tog tre resor."
		-- Joan of Arc

%
QOTD:"Vem? Mig? Nej, nej, nej !! Men jag säljer mattor."
		-- Joan of Arc

%
QOTD:"Skulle det inte vara underbart om det verkliga livet stöds kontroll-Z?"
		-- Joan of Arc

%
QOTD:"Du vill att jag ska sätta * hål * i mina öron och hänga saker från dem?Hur ... tribal. "
		-- Joan of Arc

%
QOTD:"Du är så dum att du inte ens har visdomständer."
		-- Joan of Arc

%
QOTD:Allt jag vill ha är en lite mer än jag någonsin kommer att få.
		-- Joan of Arc

%
QOTD:Allt jag vill ha är mer än min beskärda del.
		-- Joan of Arc

%
QOTD:	Blixt! Blixt! Jag älskar dig! ... Men vi bara har fjorton timmar till	rädda jorden!
		-- Joan of Arc

%
QOTD:Hur kan jag sakna dig om du inte kommer att försvinna?
		-- Joan of Arc

%
QOTD:Jag tittade ut mitt fönster och såg Kyle Pettys "bil upp och ner,då tänkte jag "En av oss är i verkliga problem.
		-- Davey Allison, on a 150 m.p.h. crash

%
QOTD:Jag älskar din outfit, kommer det i din storlek?
		-- Davey Allison, on a 150 m.p.h. crash

%
QOTD:Jag öppnade Pandoras ask, låta katten ur påsen och sättabollen på deras planhalva.
		-- Hon. J. Hacker (The Ministry of Administrative Affairs)

%
QOTD:Jag är inte en nerd - Jag är "socialt utmanade".
		-- Hon. J. Hacker (The Ministry of Administrative Affairs)

%
QOTD:Jag är inte skallig - Jag är "hår utmanade".[Jag trodde det var "annorlunda haired". Ed.]
		-- Hon. J. Hacker (The Ministry of Administrative Affairs)

%
QOTD:Jag har hört talas om civilingenjörer, men jag har aldrig träffat en.
		-- Hon. J. Hacker (The Ministry of Administrative Affairs)

%
QOTD:Om det är för högt, du är för gammal.
		-- Hon. J. Hacker (The Ministry of Administrative Affairs)

%
QOTD:Om du letar efter problem, kan jag erbjuda dig ett stort utbud.
		-- Hon. J. Hacker (The Ministry of Administrative Affairs)

%
QOTD:Ludwig Boltzmann, som tillbringar en stor del av sitt liv åt att studera statistiskmekaniker dog 1906 av hans egen hand. Paul Ehrenfest, bärandepå arbetet, dog på samma sätt 1933. Nu är det vår tur.
		-- Goodstein, States of Matter

%
QOTD:Pengar är inte allt, men åtminstone det håller barnen kontakten.
		-- Goodstein, States of Matter

%
QOTD:Min mor var resebyrån för skuld resor.
		-- Goodstein, States of Matter

%
QOTD:På en skala från 1 till 10 skulle jag säga ... oh, någonstans där inne.
		-- Goodstein, States of Matter

%
QOTD:Heliga kor gör stora hamburgare.
		-- Goodstein, States of Matter

%
QOTD:Tystnad är den enda kraft som han har lämnat.
		-- Goodstein, States of Matter

%
QOTD:Vissa människor har en av dessa dagar. Jag har haft en av dessa liv.
		-- Goodstein, States of Matter

%
QOTD:Talang gör vad den kan, geni vad det måste.Jag gör vad jag får betalt för att göra.
		-- Goodstein, States of Matter

%
QOTD:Snacka om villiga människor ... över hälften av dem är villiga att arbetaoch de andra är mer än villiga att titta på dem.
		-- Goodstein, States of Matter

%
QOTD:Skogen kan vara tyst, men det betyder inte attormarna har försvunnit.
		-- Goodstein, States of Matter

%
QOTD:Det enda enkla sättet att berätta en hamster från en gerbil är attgerbil har mer mörkt kött.
		-- Goodstein, States of Matter

%
QOTD:Du vet hur s'm människor behandlar th'r kropp som ett tempel?Tja, jag behandlar min vilja 'n KULTUR PARK ... S'great ...
		-- Goodstein, States of Matter

%
Kvalitetskontroll, n .:Säkerställa att kvaliteten på en produkt inte urartaroch lägga till kostnaden för dess tillverkning eller utformning.
		-- Goodstein, States of Matter

%
Kvalitetskontroll, n .:Processen med att testa en av 1000 enheter kommer utanfören produktionslinje för att se till att åtminstone en av 100 verk.
		-- Goodstein, States of Matter

%
kvark:Ljudet görs av en väluppfostrad anka.
		-- Goodstein, States of Matter

%
Quigley lag:Den som har någon makt över dig, oavsett hur liten, kommeratttempt att använda den.
		-- Goodstein, States of Matter

%
QWERT (kwirt) n. [MW <OW qwertyuiop, en trettonde] 1. en viktenhetlika med 13 poiuyt avoirdupois (eller 1.69 kiloliks), som vanligen används ibyggteknik 2. [Colloq.] 1/13 den belastning som en heltodlas sligo kan bära. 3. [Anat.] En smärtsam irritation i dermisi området för anus 4. [Slang] person som exciterar det i andrasymtom på en qwert.
		-- Webster's Middle World Dictionary, 4th ed.

%
Ralph Observation:Det är ett misstag att låta någon mekanisk objekt inser att duhar bråttom.
		-- Webster's Middle World Dictionary, 4th ed.

%
Slumpmässigt, N .:Liksom i antal, förutsägbart. Som i minnesaccess, oförutsägbar.
		-- Webster's Middle World Dictionary, 4th ed.

%
Ray Rule of Precision:Mät med en mikrometer. Markera med krita. Skär med en yxa.
		-- Webster's Middle World Dictionary, 4th ed.

%
Re: Grafik:En bild säger mer 10K ord - men endast de att beskriva	bilden. Knappast några uppsättningar 10K ord kan vara ett adekvatbeskrivas med bilder.
		-- Webster's Middle World Dictionary, 4th ed.

%
Realtid, adj .:Här och nu, i motsats till falska tid, som bara förekommer där och då.
		-- Webster's Middle World Dictionary, 4th ed.

%
Verkliga världen, n .:1. I programmerings, dessa institutioner där programmering kananvändas i samma mening som FORTRAN, COBOL, RPG, IBM, etc. 2. Tillprogrammerare, platsen för icke-programmerare och aktiviteter som inte har sambandprogrammering. 3. Ett universum där standard klänning är skjorta ochslips och i vilken en persons arbetstid definieras som 9 till 5. 4.Placeringen av status quo. 5. någonstans utanför ett universitet."Dålig karl, han lämnade MIT och gått in i den riktiga världen." Begagnadenedsättande av dem inte bosatt där. I samtal, samtalav någon som har skrivit den verkliga världen är inte olikt att tala om enavliden person.
		-- Webster's Middle World Dictionary, 4th ed.

%
Omvärdering, n .:En plötslig förändring i sinnet efter att ha fått reda på.
		-- Webster's Middle World Dictionary, 4th ed.

%
Receptionen, n .:Skärselden där kontors besökare är dömda att spenderaotaliga timmar läsning hundöron tillbaka frågor rörande handeltidningar som Modern Plastics, Chain Saw åldern och kyckling World,medan receptionist läser glatt sin egen branschtidningen -Kosmopolitiska.
		-- Webster's Middle World Dictionary, 4th ed.

%
Rekursion N .:Se rekursion.
		-- Random Shack Data Processing Dictionary

%
Reformeras, n .:En synagoga som stänger för det judiska helgdagar.
		-- Random Shack Data Processing Dictionary

%
Regressionsanalys:Matematiska metoder för att försöka förstå varför saker och ting är	blir värre.
		-- Random Shack Data Processing Dictionary

%
Reichel lag:En kropp på semester tenderar att förbli på semester inte påverkas aven yttre kraft.
		-- Random Shack Data Processing Dictionary

%
Reisner härskar av begrepps Inertia:Om du tror tillräckligt stor, kommer du aldrig att göra det.
		-- Random Shack Data Processing Dictionary

%
Tillförlitlig källa, n .:Killen du just träffat.
		-- Random Shack Data Processing Dictionary

%
Renning Maxim:Människan är den högsta djuret. Man gör klassificerings.
		-- Random Shack Data Processing Dictionary

%
Reporter, n .:En författare som gissar sig fram till sanningen och skingrar det med enstorm av ord.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Rykte, adj .:Vad andra inte tänker på dig.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Forskning, n .:Överväga Columbus:Han visste inte var han var på väg.När han kom dit han inte visste var han var.När han kom tillbaka han inte visste var han hade varit.Och han gjorde det på någon annans pengar.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Ansvar:Alla säger att det är ett stort ansvar som har makt. Detta ären hel del säng. Ansvaret är när någon kan klandra dig om någotgår fel. När du har makt du är omgiven av människor vars jobb detär att ta på sig skulden för dina misstag. Om de är smarta, är det.
		-- Cerebus, "On Governing"

%
Revolution, n .:En form av regering utomlands.
		-- Cerebus, "On Governing"

%
Revolution, n .:I politiken, en abrupt förändring i form av vanstyre.
		-- Ambrose Bierce

%
revolutionerande, adj .:Ompaketerade.
		-- Ambrose Bierce

%
Rhode lag:När någon princip lag, grundsats, sannolikhet, händer, omständighet,eller resultat kan inte på något sätt vara direkt, indirekt, empiriskt, elleromvägar bevisat, härledd, underförstådda, antagen, inducerad, dras,uppskattad eller vetenskapligt gissat, det kommer alltid för ändamåletbekvämlighet, ändamålsenlighet, politiska fördelar, materiell vinning, ellerpersonlig komfort, eller någon kombination av de ovanstående eller ingen av deovan, ensidigt och otvetydigt antas förkunnade, ochföljs som absolut sanning att vara onekligen, universellt, oföränderligt,och oändligt så, fram till dess att det blir fördelaktigt attantar annars kanske.
		-- Ambrose Bierce

%
Ritchies Regel:(1) Allt har ett visst värde - om du använder rätt valuta.(2) färgstänk sist längre än lack.(3) Sök och ni skall finna - men se till att det var förlorat.
		-- Ambrose Bierce

%
Robot, n .:Universitets administratören.
		-- Ambrose Bierce

%
Robusthet, adj .:Aldrig behöva säga att du är ledsen.
		-- Ambrose Bierce

%
Rockys Lemma för förebyggande Innovation:Inte resultatet är kända i förväg, finansiärer kommerförkasta förslaget.
		-- Ambrose Bierce

%
Rudd Discovery:Du vet att någon senator eller kongressledamot kunde gå hem och göra$ 300.000 till $ 400.000, men de gör det inte. Varför? Eftersom de kanstanna i Washington och göra det där.
		-- Ambrose Bierce

%
Rudin lag:Om det finns ett fel sätt att göra något, de flesta människor kommergör det varje gång.Rudin andra lag:I en kris som tvingar ett val göras mellan alternativhandlings, människor tenderar att välja den värsta möjligakurs.
		-- Ambrose Bierce

%
robust, adj .:För tung att lyfta.
		-- Ambrose Bierce

%
Regel nr 1:Boss är alltid rätt.Regel # 2:Om chefen är fel, se Regel nr 1.
		-- Ambrose Bierce

%
Rule of Creative Forskning:(1) dra aldrig vad du kan kopiera.(2) kopiera aldrig vad du kan spåra.(3) spår aldrig vad du kan klippa ut och klistra ner.
		-- Ambrose Bierce

%
Rule of Defactualization:Information försämras uppåt genom byråkratier.
		-- Ambrose Bierce

%
Rule of Feline frustration:När din katt har somnat i knät och ser fullständigtinnehåll och bedårande, kommer du plötsligt att gå tillbadrum.
		-- Ambrose Bierce

%
Rule of the Great:När människor du beundrar verkar tänka djuptankar, de förmodligen tänker lunch.
		-- Ambrose Bierce

%
Regler för Academic Deans:(1) Hide !!!!(2) Om de hittar dig, lie !!!!
		-- Father Damian C. Fandal

%
Regler för körning i New York:(1) Allt gjort medan tutande din horn är lagligt.(2) Du kan parkera var som helst om du förvandla dina fyrvägs blinkers på.(3) Ett rött ljus innebär de kommande sex bilar kan gå igenomkorsning.
		-- Father Damian C. Fandal

%
Regler för författare:Undvika run-på meningar som de är svåra att läsa. Använd inte någon dubbelnegativ. Använd semikolon korrekt, alltid använda den när det är lämpligt,och aldrig var det inte. Reserverar apostrof för det är korrekt användning ochutelämna det när det inte behövs. Inga meningsfragment. Undvik kommatecken, som äronödig. Undfly dialekt, Oberoende. Och inte börja en mening meden konjunktion. Avstava mellan SY-llables och undvika onödiga bindestreck.Skriv alla adverbiella former korrekt. Använd inte sammandragningar i formell skrift.Skriver noggrant, måste dinglande participles undvikas. Det åliggeross att undvika arkaismer. Undvika felaktiga former av verb som harsmet i språket. Aldrig, aldrig använda repetitiva uppsägningar. Om jag harberättade dig en gång, har jag sagt tusen gånger, motstå överdrift. Också,undvika besvärliga eller påverkas allitteration. Inte sträng alltför många prepositionalfraser tillsammans om du vandrar genom dalen i skuggan avdöd. "Undvik överanvändning av" citat "märken." ' "
		-- Father Damian C. Fandal

%
Runes regel:Om du inte bryr var du är, är du inte förlorat.
		-- Father Damian C. Fandal

%
Ryans lag:Gör tre korrekta gissningar följdoch du kommer att etablera dig som en expert.
		-- Father Damian C. Fandal

%
Sacher Observations:Vissa människor växer med ansvar - andra bara sväller.
		-- Father Damian C. Fandal

%
Satellit Safety Tips # 14:Om du ser en ljus strimma på himlen kommer på dig, anka.
		-- Father Damian C. Fandal

%
Sattinger lag:Det fungerar bättre om du ansluter den.
		-- Father Damian C. Fandal

%
Savage lag lämplighets:Du vill ha det dåligt, får du det dåligt.
		-- Father Damian C. Fandal

%
scenario, n .:En tänkt sekvens av händelser som ger det sammanhang isom ett affärsbeslut fattas. Scenarier kommer alltiduppsättningar av tre: bästa fall värsta fall, och i fall.
		-- Father Damian C. Fandal

%
Schapiro förklaring:Gräset är alltid grönare på andra sidan - men det äreftersom de använder mer gödsel.
		-- Father Damian C. Fandal

%
Schlattwhapper, n .:Fönstret nyans som låter sig dras ner,tvekar en sekund, snäpper sedan upp i ansiktet.
		-- Rich Hall, "Sniglets"

%
Schmidts Observation:Allt annat lika, en fet person använder mer tvålän en tunn person.
		-- Rich Hall, "Sniglets"

%
Scotts första lag:Oavsett vad som går fel, kommer det förmodligen ser rätt.Scotts andra lag:När ett fel har upptäckts och korrigerats, kommer det finnasha varit fel i första hand.Naturlig följd:Efter korrigeringen har påträffats i fel, kommer det att varaomöjligt att passa den ursprungliga kvantiteten tillbaka in iekvation.
		-- Rich Hall, "Sniglets"

%
scribline, n .:Den tomt område på baksidan av kreditkort där en underskrift går.
		-- "Sniglets", Rich Hall & Friends

%
Andra lag för taxi:Om det finns två möjliga sätt att stava en persons namn, duhämtar fel.Naturlig följd:Om det bara finns ett sätt att stava ett namn,du kommer att stava det fel i alla fall.
		-- "Sniglets", Rich Hall & Friends

%
Andra lag slutprov:I din tuffaste final - för första gången hela året - den mestdistractingly attraktiv elev i klassen kommer att sitta bredvid dig.
		-- "Sniglets", Rich Hall & Friends

%
Sekreterare hämnd:Arkivering nästan allt under "den".
		-- "Sniglets", Rich Hall & Friends

%
Seleznick teori av Holistisk medicin:Ice Cream botar alla sjukdomar. Tillfälligt.
		-- "Sniglets", Rich Hall & Friends

%
Självtest för Paranoia:Du vet att du har det när du inte kan komma på något som ärditt eget fel.
		-- "Sniglets", Rich Hall & Friends

%
Senat, n .:En kropp av äldre herrar laddade med höga tullar och förseelser.
		-- Ambrose Bierce

%
senilitet, n .:Sinnestillstånd av äldre personer med vilka man råkar oense.
		-- Ambrose Bierce

%
serendipity, n .:Den process genom vilken mänsklig kunskap är avancerad.
		-- Ambrose Bierce

%
Serocki s Striktur:Äktenskapet är alltid en kandidat sista alternativet.
		-- Ambrose Bierce

%
Shannons Observation:Ingenting är så frustrerande som en dålig situation som börjarförbättras.
		-- Ambrose Bierce

%
aktie, n .:Att ge efter, uthärda förödmjukelse.
		-- Ambrose Bierce

%
Shaws Princip:Bygga ett system som även en dåre kan använda, och endast en dåre kommervill använda den.
		-- Ambrose Bierce

%
Shedenhelm lag:Alla spår har fler stigningar än de har downhill sektioner.
		-- Ambrose Bierce

%
Shick lag:Det är inga problem en bra mirakel kan inte lösa.
		-- Ambrose Bierce

%
Silverman lag:Om Murphys lag kan gå fel, kommer det.
		-- Ambrose Bierce

%
Simon lag:Allt tillsammans faller sönder förr eller senare.
		-- Ambrose Bierce

%
Skinners Constant (eller Flannagan s Finagling Factor):Denna kvantitet som när multiplicerat med dividerat med, läggas till,eller subtraheras från svaret du fick, ger dig svaret duborde ha fått.
		-- Ambrose Bierce

%
Slick s tre lagarna av universum:(1) Ingenting i det kända universum färdas snabbare än en dålig kontroll.(2) En fjärdedel uns av choklad = fyra pounds av fett.(3) Det finns två typer av smuts: den mörka slag, vilket ärattraherad av lätta föremål, och ljuset slag, vilket ärattraheras till mörka objekt.
		-- Ambrose Bierce

%
Slous påstående:Om du gör ett jobb alltför väl, kommer du fastnar med den.
		-- Ambrose Bierce

%
Slurm, n .:Slem som samlas på undersidan av en tvål närdet sitter i skålen för länge.
		-- Rich Hall, "Sniglets"

%
Snacktrek, n ​​.:Den säregna vana, när du söker efter ett mellanmål, ständigtåtervänder till kylskåpet i hopp om att något nytt kommer att haförverkligats.
		-- Rich Hall, "Sniglets"

%
galleriets repliker:Vad skulle du säga om du hade en chans.
		-- Rich Hall, "Sniglets"

%
Sodd andra lag:Förr eller senare, är den värsta möjliga mängd omständigheteratt dyka.
		-- Rich Hall, "Sniglets"

%
Programvara, N .:Formell kväll klädsel för kvinnliga datoranalytiker.
		-- Rich Hall, "Sniglets"

%
Några punkter att komma ihåg [om djur]:(1) Gå inte att sova under stora djur, exempelvis elefanter, rhinoceri,hippopotamuses;(2) Placera inte djur med vassa tänder eller giftiga huggtänder nerframför dina kläder;(3) inte klappa vissa djur, t.ex. krokodiler och skorpioner eller hundardu just har sparkas.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
spagmumps, n .:Vilken som helst av de miljontals Styrofoam tussar som följer postorder poster.
		-- "Sniglets", Rich Hall & Friends

%
Speer 1st lag Korrekturläsning:Synligheten för ett fel är omvänt proportionell mot denantalet gånger du har tittat på det.
		-- "Sniglets", Rich Hall & Friends

%
Spence förmaning:Aldrig stuva undan på en kamikaze plan.
		-- "Sniglets", Rich Hall & Friends

%
Spirtle, n .:Den fina ström från en grapefrukt som alltid landar rätt i ögat.
		-- Sniglets, "Rich Hall & Friends"

%
Make, n .:Någon som kommer att stå dig genom alla problem duskulle inte ha haft om du hade stannat singel.
		-- Sniglets, "Rich Hall & Friends"

%
squatcho, n .:På knappen på toppen av en keps.
		-- "Sniglets", Rich Hall & Friends

%
standarder, n .:De principer som vi använder för att förkasta andras kod.
		-- "Sniglets", Rich Hall & Friends

%
statistik, n .:Ett system för att uttrycka dina politiska fördomar i övertygandevetenskaplig skepnad.
		-- "Sniglets", Rich Hall & Friends

%
Steckel härskar till framgång:Bra nog är aldrig bra nog.
		-- "Sniglets", Rich Hall & Friends

%
Steele lag:Det finns uppgifter som inte kan utföras av mer än tio mäneller färre än hundra.
		-- "Sniglets", Rich Hall & Friends

%
Steeles Plagiat av Någon filosofi:Alla ska tro på något - jag tror jag kommer att haen annan dryck.
		-- "Sniglets", Rich Hall & Friends

%
Steinbach riktlinje för Systemprogrammering:testar aldrig för ett fel som du inte vet hur man ska hantera.
		-- "Sniglets", Rich Hall & Friends

%
Stenderup lag:Ju tidigare du halkar efter, desto mer tid du har att komma ikapp.
		-- "Sniglets", Rich Hall & Friends

%
Beståndets Observation:Du behöver inte förr få huvudet ovanför vattenytan, men vad någon drardina simfötter off.
		-- "Sniglets", Rich Hall & Friends

%
Sten lag:En mans "enkla" är en annan mans "va?"
		-- "Sniglets", Rich Hall & Friends

%
strategi, n .:En omfattande plan för passivitet.
		-- "Sniglets", Rich Hall & Friends

%
Strategi:En långsiktig plan vars meriter inte kan utvärderas förrän någon gångefter de som skapar det ha lämnat organisationen.
		-- "Sniglets", Rich Hall & Friends

%
Stult rapport:Våra problem är mestadels bakom oss. Vad vi måste göra nu ärbekämpa lösningar.
		-- "Sniglets", Rich Hall & Friends

%
Dum, n .:Att förlora $ 25 på spelet och $ 25 om omedelbar uppspelning.
		-- "Sniglets", Rich Hall & Friends

%
Stör lag:90% av allt är crud.
		-- "Sniglets", Rich Hall & Friends

%
socker pappa, n .:En man som har råd att höja cain.
		-- "Sniglets", Rich Hall & Friends

%
SUN Microsystems:Nätverket är belastningen Average.
		-- "Sniglets", Rich Hall & Friends

%
solnedgång, n .:Uttalad atmosfärisk spridning av kortare våglängder,vilket resulterar i selektiv överföring under 650 nanometer medgradvis minska sol höjd.
		-- "Sniglets", Rich Hall & Friends

%
sushi, n .:När det-som-kan-still-be-alive läggs ovanpå ris ochfastspänd på med eltejp.
		-- "Sniglets", Rich Hall & Friends

%
Sushido, n .:Sättet att tonfisk.
		-- "Sniglets", Rich Hall & Friends

%
Swahili, n .:Det språk som används av National Enquirer att skriva ut sina indragningar.
		-- Johnny Hart

%
Tröja, n .:Ett plagg som bärs av ett barn när dess mamma känns kyligt.
		-- Johnny Hart

%
Swipple s Rule of Order:Den som ropar högst har ordet.
		-- Johnny Hart

%
systemoberoende, adj .:Fungerar lika dåligt på alla system.
		-- Johnny Hart

%
T-shirt av dagen:Chef för bergenUppföljning T-shirt av dagen (på samma natursköna bakgrund):Om du gillade bergen, chef för Busch!
		-- courtesy someone else

%
T-shirt av dagen:Jag är personen din mamma varnade dig omkring.
		-- courtesy someone else

%
T-shirt:Livet är * inte * en Cabaret, och sluta kalla mig kompis!
		-- courtesy someone else

%
Takt, n .:Den osagt del av vad du tänker.
		-- courtesy someone else

%
vidta kraftfulla åtgärder:Gör något som borde ha gjorts för länge sedan.
		-- courtesy someone else

%
skattekontoret, n .:Den av orättvisa.
		-- courtesy someone else

%
Skatter, n .:Av livets två visshet, den enda som kan du fåen förlängning.
		-- courtesy someone else

%
konservator, n .:En man som monterar djur.
		-- courtesy someone else

%
TCP / IP-Slang Ordlista, # 1:Gong, n: Medeltida term för dass, eller vad pased för dem på den tiden.Idag används whimsically att beskriva efterdyningarna av en bogon attack. Trori vårt samhälle som Galapagos av det engelska språket."Vogons kan läsa dig dålig poesi, men bogons gör du studerar föråldrade RFC."
		-- Dave Mills

%
lagarbete, n .:Efter att ha någon att skylla.
		-- Dave Mills

%
Technicality, n .:I en engelsk domstol en man vid namn Hem prövades för förtal att haanklagade en granne för mord. Hans exakta ord var: "Sir Thomas Holthar tagit sig en köttyxa och drabbade hans kock på huvudet, så att ensidan av hans huvud föll på ena axeln och den andra sidan på denandra axeln. "Svaranden frikändes av instruktion fördomstol, de lärda domarna anse att orden inte ut mord,för de inte bekräfta död kocken, som är bara enslutledning.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Telefon, n .:En uppfinning av djävulen som upphäver några av fördelarnaatt göra en oangenäm person hålla sitt avstånd.
		-- Ambrose Bierce

%
telepression, n .:Den djupa skuld som härrör från att veta att du inte försökertillräckligt hårt för att slå upp numret på egen hand och i stället sättabörda på katalogen assistent.
		-- "Sniglets", Rich Hall & Friends

%
Germansk:Inte nog gin.
		-- "Sniglets", Rich Hall & Friends

%
Den 357,73 Teori:Revisorer alltid avvisar räkningarmed en nedersta raden delbart med fem.
		-- "Sniglets", Rich Hall & Friends

%
Den Abrams 'Princip:Det kortaste avståndet mellan två punkter är off the wall.
		-- "Sniglets", Rich Hall & Friends

%
Den antika läran om Mind Over Matter:Jag har inget emot ... och du inte spelar någon roll.
		-- As revealed to reporter G. Rivera by Swami Havabanana

%
Skalbaggarna:Paul McCartney gamla back-up band.
		-- As revealed to reporter G. Rivera by Swami Havabanana

%
Briggs-Chase lag Program Development:För att avgöra hur lång tid det tar att skriva och felsöka enprogram, ta din bästa uppskattning, multiplicera det med två, läggen, och konvertera till nästa högre enheter.
		-- As revealed to reporter G. Rivera by Swami Havabanana

%
Konsulten förbannelse:När kunden har slagit på dig tillräckligt länge, ge honomvad han ber om, i stället för vad han behöver. Detta är mycket starkmedicin, och normalt krävs endast en gång.
		-- As revealed to reporter G. Rivera by Swami Havabanana

%
Distinktionen mellan judiska och goyish kan vara ganska subtil, somföljande citat från Lenny Bruce illustrerar:"Jag är jude. Count Basie judiska. Ray Charles är judisk.Eddie Cantors goyish. B'nai Brith är goyish. Hadassah ärJudisk. Marine Corps - tung goyish, farlig."Kool-Aid är goyish. Alla Drakes Kakor är goyish.Pumpernickel är judisk och som ni vet, är mycket goyish vitt bröd.Omedelbar potatis - goyish. Körsbär soda är mycket judisk.Mandelbiskvier är ____ mycket judisk. Fruktsallad är judisk. Lime Jell-O ärgoyish. Lime soda är ____ väldigt goyish. Släpvagn parker är så goyish attJudar inte gå nära dem ... "
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Femte regeln:Du har tagit dig alltför allvarligt.
		-- Arthur Naiman, "Every Goy's Guide to Yiddish"

%
Den första regeln för programoptimering:Gör det inte.Den andra regeln för Program Optimization (endast experter!):Gör det inte ännu.
		-- Michael Jackson

%
De fem regler för socialismen:(1) Tro inte.(2) Om du tror, ​​inte talar.(3) Om du tänker och talar, inte skriva.(4) Om du tror att tala och skriva, inte underteckna.(5) Om du tror att tala, skriva och underteckna inte bli förvånad.
		-- being told in Poland, 1987

%
Följande inordna alla fysiska och mänskliga lagar:(1) Du kan inte trycka på en sträng.(2) är inte inga fria luncher.(3) Dem som har blir.(4) Du kan inte vinna dem alla, men du säker på som fan kan förlora dem alla.
		-- being told in Poland, 1987

%
Den gyllene regeln of Arts and Sciences:Han som har guldet gör reglerna.
		-- being told in Poland, 1987

%
Den gordiska Maxim:Om en sträng har en ände, har den en annan.
		-- being told in Poland, 1987

%
Den stora Bald Swamp Hedgehog:Den stora Bald Swamp Hedgehog av Billericay displayer, i uppvaktning,hans enda tagg och gör intryck av Holiday Inn desk.Eftersom detta innebär honom stående orörlig för enorma perioderNär han är ofta äts i full skärm av The Great Bald SwampHedgehog Eater.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Heineken osäkerhetsprincip:Du kan aldrig vara säker på hur många öl du hade i går kväll.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Historien om krigföring på liknande sätt delas, även här fasernaär Retribution, Förväntan, och diplomati. Således:Vedergällning:Jag ska döda dig eftersom du dödade min bror.Förväntan:Jag ska döda dig eftersom jag dödade din bror.Diplomati:Jag kommer att döda min bror och sedan döda dig påförevändning att din bror gjorde det.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Illiterati Programus Canto 1:Ett program är väldigt lik en näsa: Ibland körs ochibland blåser.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Kennedy Constant:Inte arg - få ännu.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Lagen om brevet:Det bästa sättet att inspirera färska tankar är att försegla kuvertet.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Marinkåren:De få, stolt, de döda på stranden.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Marinkåren:De få, stolt, det inte mycket ljus.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den Modelski kedjeregeln:(1) Se intensivt på problemet i flera minuter. kliar dinhuvud vid 20-30 sekunders intervall. Försök att lösa problemet på egenHewlett-Packard.(2) Om detta titta runt på klassen. Välj en särskiltljusa utseende individ.(3) Procure en stor kedja.(4) Gå över till den valda eleven och hotar att slå honom hårtmed kedjan om han inte ger dig svaret på problemet.I allmänhet kommer han. Det kan också vara en bra idé att ge honom ett ljudstryk ändå, bara för att visa att du menar allvar.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den farligaste organisationen i Amerika idag är:(A) KKK(B) Den amerikanska nazistpartiet(C) Delta Frequent Flyer Club
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den officiella MBA handbok om visitkort:Undvik alltför pretentiösa titlar som "Lord of the Realm,Trons försvarare, Emperor of India "eller" Director of CorporatePlanering. "
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den officiella MBA handbok om att göra företagets verksamhet på ett flygplan:Fungerar inte öppet på topphemliga företag kostnads ​​dokument såvidadu tidigare har konstaterat att passageraren bredvid digär blind, en musiker på humörlindrande läkemedel, ellerolyckligt innehavaren av 1/47 kromosomen.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den officiella MBA handbok om användningen av sollampor:Använd en sollampa bara på helgerna. På så sätt, om kontoret klok killeanmärker på det plötsliga uppdykandet av din solbränna, kan du tillverkanågon historia om en sol-strök helg på någon ö Shangri-Lagillar Caneel Bay. Ingenting är mer transparent än lämnarkontor vid 11:45 på en tisdag natt, bara för att återvända en Aztec solgud vid 08:15 nästa morgon.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
The Phone Booth regel:En ensam dime blir alltid antalet nästan rätt.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den qotc (citat av con) var Liz:"Min hjärna söks ut till min lever."
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den verkliga mannens Bloody Mary:Ingredienser: vodka, tomatjuice, Tobasco, Worcestershiresås, A-1 stek sås, is, salt, peppar, selleri.Fyll en stor tumlare med vodka.Kasta alla andra ingredienser bort.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den romerska regeln:Den som säger att det inte kan göras bör aldrig avbrytaen som gör det.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Reglerna:(1) Du skall inte tillbe andra datorsystem.(2) Du skall inte uppträda Liberace eller äta vattenmelon medansitter på konsolen tangentbord.(3) Du skall inte slå användare i ansiktet, eller häftklammer deras fånigasmå kortlekar tillsammans.(4) Du skall inte bli fysiskt involverad i datorsystemet,speciellt om du redan är gift.(5) Du skall inte använda magnetband som frisbees, eller använd en skivapack som en pall för att nå en annan disk pack.(6) Du skall inte stirra på blinkande lampor för mer än enåtta timmars skift.(7) Du skall inte tala om användare som du av misstag förstörde derasfiler / backup bara för att se utseendet på sina små ansikten.(8) Du skall inte njuta avbryta ett jobb.(9) Du skall inte visa skjutvapen i datasalen.(10) Du skall inte tryckknappar "bara för att se vad som händer".
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Den termodynamikens andra lag:Om du tror att saker och ting är i en enda röra nu, vänta bara!
		-- Jim Warner

%
Den sjunde budorden för tekniker:Arbetet du inte på spänningssatt utrustning, för om vad du bör göra, din kollegaarbetare vill köpa öl för din änka och trösta henne i andrasätt.
		-- Jim Warner

%
Sjätte budet frisbee:Den största enskilda stödet till avståndet är för skivan att gå i enriktning du inte vill. (Går åt fel håll = går långt.)
		-- Dan Roddick

%
Den tredje lag Foto:Om du lyckades få några bra skott, kommer de att förstörasnär någon av misstag öppnar mörkrummet dörren och allade mörka läcker ut.
		-- Dan Roddick

%
De tre största mjukvaru lögner:(1) * Naturligtvis * ger vi dig en kopia av källan.(2) * Naturligtvis * tredjepartsleverantören vi köpte den frånkommer att fixa mikrokoden.(3) Beta testplats? Nej, * naturligtvis * du inte är en beta testplats.
		-- Dan Roddick

%
De tre Termodynamikens:(1) Du kan inte få något utan att arbeta för det.(2) Det mesta du kan åstadkomma genom att arbeta är att nollresultat.(3) Du kan endast bryta även vid absoluta nollpunkten.
		-- Dan Roddick

%
Sats: en katt har nio svansar.Bevis:Ingen katt har åtta svansar. En katt har en svans mer än ingen katt.Därför har en katt nio svansar.
		-- Dan Roddick

%
Sats: Alla positiva heltal är lika.Bevis: Tillräckligt för att visa att för varje två positiva heltal, A och B, A = B.Vidare är det tillräckligt att visa att för alla N> 0, om A och B(Positiva heltal) uppfyller (MAX (A, B) = N) då A = B.Fortsätt genom induktion:Om N = 1, då A och B, som är positiva heltal, måste båda vara en.Så A = B.Antag att satsen är sant för ett visst värde på k. Take A och B medMAX (A, B) = k + 1. Sedan MAX ((A-1), (B-1)) = k. Och följaktligen(A-1) = (B-1). Följaktligen A = B.
		-- Dan Roddick

%
Theory of Selektiv Övervakning:Den tid på dagen som du luta dig tillbaka och koppla av ären gång chefen promenader genom kontoret.
		-- Dan Roddick

%
teori, n .:System av idéer avsedda att förklara något, som valts i syfte attoriginalitet, controversialism, obegriplighet, och hur bradet kommer att se ut i tryck.
		-- Dan Roddick

%
Det finns tre sätt att få något gjort:(1) Gör det själv.(2) anlita någon att göra det åt dig.(3) Förbjud dina barn att göra det.
		-- Dan Roddick

%
De älskvärda Brits avdelning:De har också svårt att uttala `vitamin".
		-- Dan Roddick

%
Tre regler för att låta som en expert:(1) förenkling era förklaringar till den grad av värdelöshet.(2) pekar alltid ut andra ordningens effekter, men aldrig påpekanär de kan ignoreras.(3) Kom upp med tre regler för din egen.
		-- Dan Roddick

%
Timjan lag:Allt går fel på en gång.
		-- Dan Roddick

%
tidsdelning, n:En tillgång metod varigenom en dator missbruk många människor.
		-- Dan Roddick

%
Dagens Tips:Stek aldrig bacon i naken.[Korrigering: alltid stek bacon i naken; Du lär inte bränna den]
		-- Dan Roddick

%
TIPS för utövande:Spelkort har den övre halvan upp-och-ner för att hjälpa fuskare.Det finns ett begränsat antal skämt i universum.Sång är ett trick för att få folk att lyssna på musik längre ände skulle normalt.Det finns ingen musik i rymden.Folk kommer att betala för att titta på folk göra ljud.Allt på scenen bör vara större än i verkliga livet.
		-- Dan Roddick

%
idag, n .:En trevlig plats att besöka, men du kan inte stanna här länge.
		-- Dan Roddick

%
toalett toup "ee, n .:Alla rulltobak mattan som orsakar locket blir topp-tung, vilketskapa oändliga irritation manliga användare.
		-- Rich Hall, "Sniglets"

%
Toni lösning på en skuldfri Life:Om du måste ljuga för någon, det är deras fel.
		-- Rich Hall, "Sniglets"

%
överföring, n .:En befordran du får under förutsättning att du lämnar stan.
		-- Rich Hall, "Sniglets"

%
transparent, adj .:Att eller i samband med ett befintligt, nontangible objekt."Det är där, men du kan inte se det"virtuell, adj .:Att eller i samband med en konkret, obefintlig objekt."Jag kan se det, men det är inte det."
		-- Lady Macbeth.

%
resa, n .:Något som gör att du känner att du får någonstans.
		-- Lady Macbeth.

%
"Lita på mig":Översättning av det latinska "varning emptor."
		-- Lady Macbeth.

%
Sanningsenliga, adj .:Dum och analfabeter.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Tsort s Konstant:1.67563, eller exakt 1,237.98712567 gånger skillnaden mellanavståndet till solen och vikten av en liten orange.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
Turnaucka lag:Uppmärksamheten span av en dator är endast så länge som desselsladd.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
Tussman lag:Ingenting är så oundviklig som ett misstag vars tid har kommit.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
US A .:"Tala inte till busschauffören."Tyskland:"Det är strängt förbjudet för passagerare att tala till föraren."England:"Du uppmanas att avstå från att tala till föraren."Skottland:"Vad har du att vinna genom att tala till föraren?"Italien:"Svara inte föraren."
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
Udall fjärde lag:Alla ändringar eller reform du kommer att få konsekvenser diginte gillar.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
Uncle Eds tumregel:Använd aldrig tummen för en regel.Du kommer antingen slå den med en hammare eller få en flisa i den.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
Underliggande Principen om socio Genetics:Överlägsenhet är recessivt.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
förstå, v .:För att nå en punkt, i utredning av något ämne, vid vilkendu upphör att undersöka vad som verkligen är närvarande, och verka pågrundval av egen intern modell istället.
		-- Terry Pratchett, "The Light Fantastic" (slightly modified)

%
Orättvisa djurnamn:
		-- Gary Larson

%
illojal konkurrens, n .:Att sälja billigare än vad vi gör.
		-- Gary Larson

%
union, n .:En avgiftsbetalande klubbarbetare svinga strejkledningen.
		-- Gary Larson

%
Universum, n .:	Problemet.
		-- Gary Larson

%
University, n .:Som en programvara hus, förutom programvarans gratis, och det är användbart,och det fungerar, och om det bryter de kommer snabbt berätta hur man rättardet, och ...[Okej, okej, jag lämnar den, men jag tror att du förstörtrovärdigheten för hela förmögenhet programmet. Ed.]
		-- Gary Larson

%
Namnlösa lag:Om det händer, måste det vara möjligt.
		-- Gary Larson

%
oändlig rikedom, n .:Vad du lämnade ut den 15 april.
		-- Gary Larson

%
Användar n .:En programmerare som kommer att tro något du säga till honom.
		-- Gary Larson

%
användaren, n .:Ordet professionella datoranvändare använder när de menar "idiot".[Jag har alltid trott "datorexpert" var frasen hackare används när de betydde "idiot". Ed.]
		-- Dave Barry, "Claw Your Way to the Top"

%
semester, n .:En två veckors binge vila och avkoppling så intensiv attdet tar ytterligare 50 veckor efter återhåll workadaylivsstil att återhämta sig.
		-- Dave Barry, "Claw Your Way to the Top"

%
Vail andra Axiom:Mängden arbete som skall utföras ökar i proportion tillmängd arbete som redan utförts.
		-- Dave Barry, "Claw Your Way to the Top"

%
Van Roy lag:Ett obrytbart leksak är användbart för att bryta andra leksaker.
		-- Dave Barry, "Claw Your Way to the Top"

%
Van Roy lag:Ärlighet är den bästa politiken - det finns mindre konkurrens.Van Roy Truism:Livet är en rad omständigheter utanför din kontroll.
		-- Dave Barry, "Claw Your Way to the Top"

%
Vanilj, adj .:Vanlig smak, standard. Se SMAK. När de används av mat,mycket ofta betyder inte att maten är smaksatt med vaniljextrahera! Till exempel "vaniljsmak vann ton soppa" (eller helt enkelt"Vanilj vann ton soppa") betyder vanlig vann ton soppa, till skillnad från hotoch sura vann ton soppa.
		-- Dave Barry, "Claw Your Way to the Top"

%
Velilind lagar Experiment:(1) Om reproducerbarhet kan vara ett problem, genomföra testet endast en gång.(2) Om en rät linje passning krävs, får endast två datapunkter.
		-- Dave Barry, "Claw Your Way to the Top"

%
Viking, n .:1. våga skandinaviska sjömän, utforskare, lycksökare,entreprenörer världsberömda för sin aggressiva, nautisk importföretag, högt belånade uppköp och blå ögon.2. Blodtörstigt hav pirater som härjade norra Europa börjari den 9: e århundradet.Hagar anmärkning: Den första definitionen är mycket föredragna; den andra användsendast av missnöjda, de avundsjuka och missnöjda ägare av vattnetfast egendom.
		-- Dave Barry, "Claw Your Way to the Top"

%
VMS, n .:Världens främsta fleranvändar äventyrsspel.
		-- Dave Barry, "Claw Your Way to the Top"

%
vulkan, n .:Ett berg med hicka.
		-- Dave Barry, "Claw Your Way to the Top"

%
Salva Teori:Det är bättre att ha lobbed och förlorat än att aldrig ha lobbed alls.
		-- Dave Barry, "Claw Your Way to the Top"

%
vuja de:Känslan av att du har * aldrig *, * någonsin * varit i den här situationen tidigare.
		-- Dave Barry, "Claw Your Way to the Top"

%
Walters "Rule:Alla flygbolag flygningar avgår från grindarna mest avlägsna fråncentrala terminalen. Ingen någonsin hade en reservationpå ett plan som lämnade Gate 1.
		-- Dave Barry, "Claw Your Way to the Top"

%
Watson lag:Tillförlitligheten av maskiner är omvänt proportionell mot denantal och betydelse av alla personer som tittar på det.
		-- Dave Barry, "Claw Your Way to the Top"

%
"Vi kommer att undersöka saken"Vid tiden hjulen gör ett helt varv, viantar att du kommer att ha glömt om det också.
		-- Dave Barry, "Claw Your Way to the Top"

%
vi:Den enskilt viktigaste ordet i världen.
		-- Dave Barry, "Claw Your Way to the Top"

%
vapen, n .:Ett index på bristande utveckling av en kultur.
		-- Dave Barry, "Claw Your Way to the Top"

%
Wedding, n:En ceremoni där två personer åtar sig att bli en, åtaratt bli ingenting och ingenting förbinder sig att bli försvarbar.
		-- Ambrose Bierce

%
Weed s Axiom:frågar aldrig två frågor i ett affärsbrev.Svaret kommer att diskutera den där du ärminst intresserade och säger ingenting om den andra.
		-- Ambrose Bierce

%
Weiler lag:Ingenting är omöjligt för den som inte har att göra det själv.
		-- Ambrose Bierce

%
Weinberg första lag:Framsteg görs endast varannan fredagar.
		-- Ambrose Bierce

%
Weinberg princip:En expert är en person som undviker de små fel medansvepande till den stora vanföreställning.
		-- Ambrose Bierce

%
Weinberg andra lag:Om byggare byggde byggnader hur programmerare skrev program,då den första hackspett som kom längs skulle förstöra civilisationen.
		-- Ambrose Bierce

%
Weiner lag av bibliotek:Det finns inga svar, bara korsreferenser.
		-- Ambrose Bierce

%
välanpassade, adj .:Förmågan att spela bridge eller golf som om de vore spel.
		-- Ambrose Bierce

%
Westheimer s Discovery:Ett par månader i laboratoriet kan ofta spara enpar timmar i biblioteket.
		-- Ambrose Bierce

%
När frågade definitionen av "pi":Matematikern:Pi är det tal som uttrycker förhållandet mellanomkretsen av en cirkel och dess diameter.Fysikern:Pi är 3.1415927, plus eller minus 0,000000005.Ingenjören:Pi är omkring 3.
		-- Ambrose Bierce

%
Whistler lag:Du vet aldrig vem som har rätt, men du alltid veta vem som är ansvarig.
		-- Ambrose Bierce

%
Vit uttalande:Tappa inte modet!Owens Kommentar till Whites uttalande:... De kanske vill klippa ut ...Byrds Tillägg till Owens Kommentar:... Och de vill undvika en lång sökning.
		-- Ambrose Bierce

%
Whitehead lag:Det självklara svaret är alltid förbises.
		-- Ambrose Bierce

%
Wiker lag:Regeringen expanderar för att absorbera intäkter och lite till.
		-- Ambrose Bierce

%
Wilcox lag:En klapp på axeln är bara några centimeter från en spark i byxorna.
		-- Ambrose Bierce

%
William Safire arbetsordning för författare:Kom ihåg att aldrig dela en infinitiv. Den passiva röst ska aldrig varaBegagnade. Placera inte uttalanden i negativ form. Verb måste hålla medsina undersåtar. Korrekturläsa noga för att se om du ord ut. Om du läsaditt arbete, kan du hitta på rereading en hel del upprepningar kan varaundvikas genom rereading och redigering. En författare får inte flytta din synpunktse. Och inte börja en mening med en konjunktion. (Kom också ihåg enpreposition är ett fruktansvärt ord för att avsluta en mening med.) Inte överutropstecken !! Placera pronomen så nära som möjligt, särskilt i de långameningar, per 10 eller fler ord till sina föregångare. Skriver noga,dinglande participles måste undvikas. Om ett ord är olämpligt i slutet aven mening, är en länk verb. Ta tjuren vid handen och undvika att blandametaforer. Undvik trendiga talesätt som låter flagnande. Alla ska varanoga med att använda en enda pronomen med singular substantiv i sitt skrivande.plocka alltid på rätt idiom. Adverbet följer alltid verbet. Sistamen inte minst, undvika klichéer som pesten; söka livskraftiga alternativ.
		-- Ambrose Bierce

%
Williams och Holland lag:Om tillräckligt med uppgifter samlas in, kan något bevisas av statistiskmetoder.
		-- Ambrose Bierce

%
Wilner Observations:Alla samtal med en potatis bör ske i privat.
		-- Ambrose Bierce

%
Wit, n .:Saltet med vilken den amerikanska Humorist skämd sin matlagnings... Genom att lämna ut det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
wok, n .:Något att thwow på wabbit.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
wolf, n .:En man som känner till alla anklarna.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Wombat lagar Dataval:(1) Om det inte körs Unix, glöm det.(2) Alla datorer designen över 10 år gammal är föråldrad.(3) Allt som IBM är skräp. (Se nummer 2)(4) Den minsta acceptabla processorkraft för en enskild användare är enVAX / 780 med en flyttalsaccelerator.(5) Alla datorer med en mus är värdelös.
		-- Rich Kulawiec

%
Woodwards lag:En teori är bättre än dess förklaring.
		-- Rich Kulawiec

%
Woolsey-Swanson Regel:Folk skulle hellre leva med ett problem som de inte kanlösa snarare än att acceptera en lösning de kan inte förstå.
		-- Rich Kulawiec

%
Arbete Regel: tjänstledighet (för en operation):Vi har slutat tillåter denna praxis. Vi vill avskräcka någontankar som du kanske inte behöver alla vad du har, och du bör inteöverväga att ha något tas bort. Vi anställde dig som du är, och att hanågot bort skulle säkert göra dig mindre än vi räknat med.
		-- Rich Kulawiec

%
arbete, n .:Den välsignade respit från skrikande barn ochsåpoperor som du faktiskt få betalt.
		-- Rich Kulawiec

%
Värsta månad 1981 för utförsåkning:Augusti. Hissen linjer är den kortaste, men.
		-- Steve Rubenstein

%
Värsta månaden på året:Februari. Februari har bara 28 dagar i det, vilket innebär att omdu hyr en lägenhet, betalar du för tre hela dagar duinte får. Försök att undvika Februarys när det är möjligt.
		-- Steve Rubenstein

%
Värsta svar på en kris, 1985:Från en läsare "Q och en kolumn i TV Guide:" Om vi ​​engagerai ett kärnvapenkrig skulle elektromagnetiska pulser från exploderande bomberskada mina videoband? "
		-- Steve Rubenstein

%
Värsta Vegetabiliska of the Year:De brysselkål. Detta är också den värsta vegetabiliska nästa år.
		-- Steve Rubenstein

%
skrivskyddsfliken, n .:Ett litet klistermärke som skapats för att täcka fula hack slarvigt kvarav skivtillverkare. Användningen av fliken skapar ett felmeddelandedå och då, men dess estetiska värde långt uppväger den momentanaolägenhet.
		-- Robb Russon

%
WYSIWYG:	Vad du ser är vad du får.
		-- Robb Russon

%
XIIdigitation, n .:Bruket att försöka bestämma året en film gjordesgenom att dechiffrera de romerska siffrorna i slutet av krediterna.
		-- Rich Hall, "Sniglets"

%
År, n .:En period av trehundrasextiofem besvikelser.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Yinkel, n .:En person som kammar sitt hår över hans kala fläck, hoppas ingenkommer att märka.
		-- Rich Hall, "Sniglets"

%
jojo, n .:Något som är tillfälligt kan upp men normalt nedåt.(Se även Computer).
		-- Rich Hall, "Sniglets"

%
Zäll s lagar:(1) Varje gång du får en munfull varm soppa, nästa sak du görkommer att vara fel.(2) hur länge en minut är, beror på vilken sida av badrummetdörr du är på.
		-- Rich Hall, "Sniglets"

%
nit, n .:Kvalitet ses i nyutexaminerade - om du är snabb.
		-- Rich Hall, "Sniglets"

%
Noll fel, n .:Resultatet av att stänga ner en produktionslinje.
		-- Rich Hall, "Sniglets"

%
Zymurgy lag av frivilligt arbete:Människor är alltid tillgängliga för arbete i förfluten tid.
		-- Rich Hall, "Sniglets"

%
Obscurism:Bruket av peppe vardagen med oklarreferenser som ett subliminalt sätt att visa upp både en utbildningoch en önskan att ta avstånd från en värld av masskultur.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
mcjob:En låg lön, låg prestige, låg-nytta, ingen framtida jobb itjänstesektor. Ofta anses vara en tillfredsställande karriär val avde som har aldrig haft en.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Fattigdom Jet Set:En grupp människor som ges till kronisk resande på bekostnad avlångsiktiga jobb stabilitet eller ett permanent uppehållstillstånd. Tenderar att ha dömtoch extremt dyra telefonsamtals relationer med människor som heterSerge eller Ilyana. Tenderar att diskutera frequent flyer program på fester.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Historisk Underdosering:Att leva i en tid när ingenting verkar hända.Större symtom beroende av tidningar, tidskrifter och TV-nyheternasändningar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Historiskt Överdosering:Att leva i en tid då alltför mycket verkar hända.Större symtom beroende av tidningar, tidskrifter och TV-nyheternasändningar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Historical slumming:Handlingen att besöka platser som diners, skorstenindustriområden, byar - platser där tiden tyckshar frysts många år tillbaka - så att uppleva lättnad nären återgår till "nuet."kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Brazilification:Den växande klyftan mellan rika och fattiga ochåtföljande försvinnande av medelklassen.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Vaccinerade Time Travel:Att fantisera om att resa bakåt i tiden, men baramed rätt vaccinationer.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Decade Blandning:I kläder: det urskillningslösa kombination av två eller fleraföremål från olika decennier för att skapa en personlig stämning: Sheila =Mary Quant örhängen (1960) + kork Wedgie plattform visar (1970) +svart skinnjacka (1950 och 1980).kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Kalvkött-gödning Pen:Små, trånga kontorsarbetsplatser byggda avtygklädd demonterbart vägg partitioner och bebos av juniorpersonal. Uppkallad efter den lilla preslaughter bås som används avboskapsindustrin.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Emotionell Ketchup Burst:Tappning av åsikter och känslor i sig såatt de explosionsartat brista ut alla på en gång, chockerande och förvirrandearbetsgivare och vänner - varav de flesta trodde det var bra.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Blödning hästsvans:En äldre, utsålda baby boomer som sörjer för hippie ellerpresellout dagar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Boomer Avund:Avund av materiell rikedom och långväga material säkerhetupplupna av äldre medlemmar av de stora åldersklasserna genomlyckliga födslar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Clique Underhåll:Behovet av en generation att se nästa led detså bristfällig så att stärka sin egen kollektiva ego: "Barn idag göraingenting. De är så apatisk. Vi brukade gå ut och protestera. Allade gör är butik och klaga. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Konsensus Terrorism:Den process som avgör tjänstgörande attityder och beteenden.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Sick Building Migration:Tendensen hos yngre arbetstagare att lämna eller undvika jobb iohälsosamma kontorsmiljöer eller arbetsplatser som berörs av de sjukaBuilding Syndrome.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Recurving:Lämnar ett jobb att ta en annan som betalar mindre men placerar entillbaka på inlärningskurvan.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Ozmosis:Oförmåga ett jobb att leva upp till en självbild.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Effekt Mist:Tendensen av hierarkier i kontorsmiljöer att diffusaoch hindra skarpa artikulation.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Overboarding:Överkompensation farhågor om framtiden genom att kastahuvudstupa in i ett jobb eller livsstil till synes orelaterade till sintidigare liv intressen: dvs Amways försäljning, aerobics, den republikanskaparti, en karriär i lag, kulter, McJobs ....kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Jordfärger:En ungdomlig grupp intresserad av vegetarianism, tie-färgadekläder, milda droger, och bra stereoutrustning. Allvarlig,ofta saknar humor.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Ethnomagnetism:Tendensen hos unga människor att leva i känslomässigtdemonstrativa, mer ohämmade etniska stadsdelar: "Du skulle inteförstå det där, mor - de * kram * där jag bor nu. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Mid-Twenties Uppdelning:En period av mental kollaps förekommer i sina tjugoårsåldern,ofta orsakas av en oförmåga att fungera utanför skolan ellerstrukturerade miljöer tillsammans med en realisering av en Essentialensamhet i världen. Ofta markerar induktion i ritualfarmaceutisk användning.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Successophobia:Rädslan att om man är framgångsrik, då ens personliga behovkommer att glömmas bort och kommer inte längre att ha sina barnsliga behovsörjt för.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Säkerhet Net-ism:Tron att det alltid kommer att vara en ekonomisk och känslomässigskyddsnät för att buffra livets ont. Vanligtvis föräldrar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Skilsmässa Antagande:En form av skyddsnät-ism, tron ​​att om ett äktenskapinte fungerar, då är det inget problem eftersom partner kan helt enkeltsöka en skilsmässa.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Anti-Sabbatical:Ett jobb tas med den enda avsikten att stanna bara för enbegränsad tidsperiod (ofta ett år). Avsikten är vanligtvis atthöja tillräckligt med pengar för att delta i en annan, mer meningsfull aktivitetsåsom akvarell skissa på Kreta, eller utforma dator stickatröjor i Hongkong. Arbetsgivarna är sällan informerade om avsikter.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Lagstadgade Nostalgia:Att tvinga en kropp av människor att ha minnen de intefaktiskt besitter: "Hur kan jag vara en del av 1960-talet generation när jaginte ens kommer ihåg något av det? "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Nu Denial:Att säga sig att den enda gången värt att leva i är det förflutna ochatt den enda gången som någonsin kan vara intressant igen är framtiden.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Bambification:Den mentala omvandling av kött och blod levande varelser iseriefigurer som har borgerliga judisk-kristna attityder ochmoral.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Sjukdomar för Kisses (Hyperkarma):En djupt rotad övertygelse om att straff på något sätt alltid kommer att varamycket större än de brott: ozonhål för nedskräpning.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Spectacularism:En fascination för extrema situationer.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
hemlöshet:En filosofi som innebär en avstämning sig med minskandeförväntningar på materiell rikedom: "Jag har gett upp att vilja göra endöda eller vara en bigshot. Jag vill bara att finna lycka och kanske öppnaupp en liten vägkanten kafé i Idaho. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Status Substitution:Använda ett objekt med intellektuell eller mode prägel tillsubstitut för ett objekt som är bara dyr "Brian, du lämnadekopia av Camus i din broders BMW. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Survivulousness:Tendensen att visualisera sig njuter av att vara den sistaperson på jorden. "Jag skulle ta en helikopter upp och kasta mikrovågsugnarner på Taco Bell. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Platonska Shadow:En icke-sexuellt vänskap med en medlem av det motsatta könet.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Mental Ground Zero:Den plats där en visualiserar sig under droppav atombomben; ofta ett köpcentrum.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Cult of Aloneness:Behovet av autonomi till varje pris, vanligtvis på bekostnad avlångsiktiga relationer. Ofta orsakas av alltför högandras förväntningar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Celebrity Schadenfreude:Lurid spänning som härrör från att tala om kändis dödsfall.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Kejsarens nya Mall:Den populära uppfattningen att köpcentra finns på insidan endastoch har ingen yttre. Upphävandet av visuella misstro alstradeav detta begrepp tillåter konsumenter att låtsas att de stora, cementblock kastats in sin omgivning inte i själva verket existerar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Poorochrondria:Hypochrondria härrör från att inte ha sjukförsäkring.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Personliga Tabu:En liten regel för att leva, som gränsar till en vidskepelse, attgör att man kan klara av vardagen i frånvaro av kulturella ellerreligiösa dictums.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Arkitektonisk matsmältningsbesvär:Den nästan tvångs behov av att leva i en "cool"arkitektoniska miljön. Ofta relaterade objekt av fetischinkluderar inramade svartvita konstfotografi (Diane Arbus afavorit); förenklat furumöbler; matt svart högteknologiska objekt sådanasom TV-apparater, stereo och telefon; låg effekt omgivande ljus; en lampa,stol eller bord som anspelar på 1950-talet; snittblommor med komplexanamn.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Japanska Minimalism:Den oftast erbjuds inredning estetiska används avrotlösa karriär-hopping ungdomar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Bröd och kretsar:Den elektroniska eran tendens att visa partipolitik som corny -inte längre är relevanta av meningsfull eller användbar för moderna samhällsfrågor,och i många fall farliga.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Väljare kvarter:Försöket är dock meningslöst, att registrera oliktänkande mednuvarande politiska systemet genom att helt enkelt inte rösta.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Armanism:Efter Giorgio Armani; en besatthet med imitera sömlösaoch (ännu viktigare) * kontrollerad * etos italienska couture. Tycka omJapanska Minimalism, Armanism speglar en djup inre behov avkontrollera.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Dålig Flytkraft:Insikten om att en var en bättre person vid en hade mindrepengar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Musikalisk hårklyverier:Handlingen att klassificera musik och musiker i patologisktPicayune kategorier: "Wien Franks är ett bra exempel på urbanvit syra fold revivalism korsas med ska. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
101-ism:Tendensen att plocka isär, ofta in i minsta detalj, allaaspekter av livet med hjälp av halv förstås pop psykologi som ett verktyg.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Yuppie Wannabes:Ett X generation grupp som tror myten om en yuppielivsstil är både tillfredsställande och livskraftiga. Tenderar att vara mycket iskuld, som deltar i någon form av missbruk, och visar en viljaatt prata om Armageddon efter tre drinkar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Ultra Short Term Nostalgia:Hemlängtan för extremt senaste tiden: "Gud, verkade sakerså mycket bättre i världen förra veckan. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Uppror Uppskjutande:Tendensen i en ungdom att undvika traditionellt ungdomligaktiviteter och konstnärliga upplevelser för att få allvarliga karriärerfarenhet. Ibland resulterar i sorg för förlorade ungdom vid caålder trettio, följt av dumma hårklippning och dyrt skämt-inducerandegarderober.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Iögonfallande Minimalism:En livsstil taktik liknar Status Byte. Denonownership av materiella varor prunkade som ett tecken på moralisk ochintellektuell överlägsenhet.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Caf 'e Minimalism:Att ansluta sig till en filosofi av minimalism utan att sättai praktiken någon av dess grundsatser.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
O'Propriation:Inkluderandet av reklam, förpackning, och underhållningjargong från tidigare epoker i dagligt tal för ironisk och / eller komiskaeffekt: "Kathleen Favorit Dead Kändisar på fest fanns massor o'fun" eller"Dave verkligen tänker på sig själv som en zany, nötig, knäpp, och våghalskille, inte han? "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Air Familj:Beskriver falsk känsla av gemenskap upplevde bland medarbetarei en kontorsmiljö.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
skruva:Obehag drabbat ungdomar från gamla människor som inte ser någonironi i deras gester. "Karen dog tusen dödsfall som hennes fargjorde en stor show av smaka en nyligen tillverkad flaska vininnan man tillåter den att hällas som familjen satt i Steak Hut.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Recreational slumming:Bruket att delta i fritidsaktiviteterav en klass man uppfattar som lägre än den egna: "Karen Donald!Låt oss gå bowling ikväll! Och oroa dig inte om skor ... tydligenkan du hyra dem. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Conversational slumming:Den självmedveten åtnjutande av en viss konversationjust för sin brist på intellektuell stringens. En stor spin-offaktivitet Recreational slumming.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Occupational slumming:Ta ett jobb väl under en skicklighet eller utbildningsnivåsom ett medel för reträtt från vuxna ansvar och / eller undvikamisslyckande i ett verkliga yrke.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Anti-Offer Enhet:En liten modetillbehör som bärs på en annarskonservativ dräkt som tillkännager för världen att man fortfarande har engnista av individualitet brinnande inuti: 1940 retro band och örhängen(På män), feministiska knappar, näsring (kvinnor), och nu nästanhelt utrotade teeny weeny "rattail" frisyr (båda könen).kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Närings slumming:Mat vars njutning beror inte från smak men från enkomplex blandning av klass konnotationer, nostalgi signaler ochförpacknings semiotik: Katie och jag köpte denna tub av Multi-Whip iställetverkliga piska grädde eftersom vi trodde petroleumdestillat piskaTaklagsfest verkade sorts mat som flygvapen fruar stationerade iPensacola tillbaka i början av sextiotalet skulle föda sina män tillfira en karriär befordran.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Tele-Parabilizing:Moral som används i vardagen som härrör från tv-serien tomter:"Det är precis som episoden där Jan förlorar sina glasögon!"kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
QFM:Quelle mode misstag. "Det var verkligen QFM. Jag menar målarebyxor? Det är 1979 obegripligt. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Me-ism:En sökning av en individ, i avsaknad av utbildning itraditionella religiösa trossatser, att formulera en skräddarsyddreligion själv. Oftast ett hopkok av reinkarnation,personlig dialog med en nebulously definierad gud siffra, naturalism,och karmiska öga för ögon attityder.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Pappers Rabies:Överkänslighet mot nedskräpning.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Bradyism:En multisibling känslighet härrör från att ha vuxit upp istora familjer. En sällsynthet i dem som är födda efter cirka 1965,symptom på Bradyism omfatta en anordning för psyk, emotionellindragning i situationer med överbeläggning, och en djupt känt behov av enväldefinierade personliga utrymme.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Svarta hål:Ett X generation grupp mest känd för sin besittningnästan helt svarta garderober.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Svarta Dens:Där svarta hål lever; ofta ouppvärmda lager med Day-Glosprutmålning, stympade skyltdockor, Elvis referenser, dussintalsfulla askkoppar, spegel skulpturer och Velvet Underground musikspelar i bakgrunden.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Strange Reproduktion:Att ha barn för att kompensera för det faktum att man inte längretror på framtiden.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Squires:Den vanligaste X generation grupp och den enda undergruppges till avel. Squires finns nästan uteslutande i par ochkänns igen på sina desperata försök att skapa ett sken avEisenhower-eran plenitude i det dagliga livet i ansiktet avorimliga bostadspriser och två lediga livsstilar. Squires tenderar att varakontinuerligt ut från deras glupskt tillgrepps strävanmöbler och prylar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Fattigdom lurar:Finansiell paranoia ingjutit i avkomma av depression-eranföräldrar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Pull-the-Plug, Skiva Pie:En fantasi där en avkomma stämmer upp mentalt dennettoförmögenhet på sina föräldrar.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Underdogging:Tendensen att nästan alltid sida med underdog i engiven situation. Konsumenten uttrycket för denna egenskap ärinköp av mindre framgångsrika, "ledsen" eller misslyckas produkter: "Jag vetDessa Wien Franks är hjärtsvikt på en pinne, men de var så tråkigttittar upp mot alla andra yuppie livsmedel som jag bara var tvungen attköp dem."kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
2 + 2 = 5-ism:Grottkrypning till en målinriktad marknadsföring strategi som syftar till sig själv efterhåller ut under en lång tidsperiod. "Åh, okej, jag ska köpa dindum cola. Nu lämnar mig ensam. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Alternativet Förlamning:Tendensen, när det ges obegränsade valmöjligheter, att ingen.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Personlighet Tithe:Ett pris som betalas för att bli ett par; tidigare underhållandemänniskor bli tråkigt: "Tack för att bjuda in oss, men Noreen och jagkommer att titta på bestick kataloger i kväll. Efteråt ska viatt titta på shoppingkanal. "kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Jack and Jill Party:A Squire tradition; baby shower som båda män ochväninnor inbjuds i motsats till endast kvinnor. fördubblatsköpkraft bisexuella närvaro ger gåva värden upp tillEisenhower-eran standarder.kultur "
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
Down-Nesting:Tendensen hos föräldrar att flytta till mindre, gästrummet fritthus efter barnen har flyttat för att undvika barn i åldern20 till 30 som har boomeranged hem.
		-- Douglas Coupland, "Generation X: Tales for an Accelerated

%
greenrd lagEvey post nedvärderande någon annans stavning eller grammatik, eller laudingen egen stavning eller grammatik, oundvikligen kommer att innehålla en stavning ellergrammatiska fel.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
intaxication:Eufori på att få en skatteåterbäring, som varar tills man inserdet var dina pengar till att börja med.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
reintarnation:Kommer tillbaka till livet som en lantis.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
bozone, n .:Ämnet som omger dumma människor som stoppar goda idéerfrån att tränga in. Den bozone skiktet olyckligtvis visar få teckenatt bryta ned inom en snar framtid.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
cashtration, n .:Handlingen att köpa ett hus, vilket gör ämnet ekonomisktimpotent på obestämd tid.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
giraffiti:Vandalism sprayat mycket, mycket hög.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
sarchasm:Klyftan mellan författaren sarkastisk kvickhet och den person sominte få det.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
inoculatte:Att ta kaffe intravenöst när du kör sent.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
hipatitis:Terminal svalka.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
osteopornosis:En degenererad sjukdom.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
Karmageddon:Det är som när alla sänder ut alla dessa verkligen dåligvibbar, eller hur? Och sedan, som, jorden exploderar och det är, enallvarlig bummer.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
decafalon, n .:Den krävande händelse av att ta sig igenom dagen förbrukar endasom är bra för dig.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
glibido:Alla samtal och ingen åtgärd.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
Dopeler effekt:Tendensen dumma idéer att verka smartare när de kommer på digsnabbt.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
arachnoleptic passform, n .:Desperata dans som utförs precis efter att du har av misstag gåttgenom ett spindelnät.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
Beelzebug, n .:Satan i form av en mygga, som hamnar i sovrummet påtre på morgonen och kan inte kastas ut.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
caterpallor, n .:Färgen du slår efter att hitta en halv grub i frukten dumat.
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
De Arrogant Worms beskriva Kanada:  Våra berg är mycket spetsiga;  våra prärier inte är det.  Resten är ganska ojämn,  men man, vi har en hel del!    - Från "Kanada är verkligen Big"
		-- greenrd in http://www.kuro5hin.org/comments/2002/4/16/61744/5230?pid=5#6

%
