100 hinkar med bitar på bussen100 hinkar med bitarTa en ner, kort det till jordFF hinkar bitar på bussenFF hinkar bitar på bussenFF hinkar bitarTa en ner, kort det till jordFE hinkar bitar på bussenoändlighet ...
		-- ``Cities in Dust'', "Tinderbox", Siouxsie & the Banshees.

%
99 block av crud på disken,99 block av crud!Du patch en bugg, och dumpa det igen:100 block av crud på skivan!100 block av crud på disken,100 block av crud!Du patch en bugg, och dumpa det igen:101 block av crud på skivan! ...
		-- ``Cities in Dust'', "Tinderbox", Siouxsie & the Banshees.

%
En bit av talkÄr alltid walcum
		-- Ogden Nash

%
En ruta utan gångjärn, nyckel, eller lock,Ändå gyllene skatt insidan dolde.
		-- J. R. R. Tolkien

%
Ett gäng pojkarna kikhosta det i Malemute saloon;Grabben som hanterar speldosa var slå en Jag-tid tune;Baksidan av stapeln, i en solospel, satt farliga Dan McGrew,Och titta på hans lycka var hans ljus o'-kärlek, damen som är känd som Lou.
		-- Robert W. Service

%
En kusin till mig sa en gång om pengar,pengar är alltid där men fickorna förändras;det är inte i samma fickorna efter en förändring,och det är allt som finns att säga om pengar.
		-- Gertrude Stein

%
En Elbereth Gilthoniel,silivren Penna m 'irielo Menel aglar elenath!Na chaered palan-d 'irielo galadhremmin ennorath,Fanuilos, le linnathonnef aear, s 'i Nef aearon!
		-- J. R. R. Tolkien

%
En montör passar; Även om syndare syndEn skär snitt; Och späd tunnaOch ett flygplan Spotter fläckar; Och pappersläskpapper blotEn barnvakt jag har aldrig ännuBaby-sitter - Hade bokstäver låtMen en utter OTs aldrig. Eller sett en utter ot.Smet fladdermöss(Eller skingrar scats);En trädgårdsskjul är för ingjutning;Men ingen har hittatEn knöl bundenEller fångas en utter Otting.
		-- Ralph Lewin

%
A är för awk, som löper som en snigel, ochB är för biff, som läser all din e-post.C är för cc, som hackare minns, medanD är för dd kommandot som gör allt.E är för emacs, som rebinds dina nycklar, ochF är för fsck, som bygger om dina träd.G är för grep, en smart detektiv, medanH är för stopp, vilket kan verka defekt.Jag är för strecksatsen som sällan roar, ochJ är för gå, som ingen använder.K är för döda, vilket gör dig till chefen, medanL är för lex, som saknas i DOS.M är för mer, varifrån en mindre var fött, ochN är för fin, som det egentligen inte.Nollan är för OD, som skriver ut saker vackert, medanP är för passwd, som läser in strängar två gånger.Q är för kvot, en Berkeley-typ fabel, ochR är för ranlib för sortering ar bord.S är för pass, som försöker förringa, medanT är för sant, som gör mycket lite.U är för uniq, som används efter sortera ochV är för VI, som är svår att avbryta.W är för whoami, som talar om ditt namn, medanX är, ja, X, av tvivelaktig berömmelse.Y är för ja, vilket gör ett intryck, ochZ är för zcat, som hanterar kompression.
		-- THE ABC'S OF UNIX

%
En dam med en av hennes öron tillämpasTill en öppen nyckelhål hört, inne,Två kvinnliga gossips i converse fri -Ämnet engagera dem var hon."Jag tror", sade en, "och min man tyckerAtt hon är en nyfikna, nyfikna minx! "Så snart inte mer av det hon kunde höraDamen, upprörd, bort hennes öra."Jag kommer inte att stanna", sade hon med en tånglake,"Att höra min karaktär ljög om!"
		-- Gopete Sherany

%
Ett litet ord av tveksamt nummer,En fiende att vila och fredlig slummer.Om du lägger till en "s" till detta,Stor är den metamorfos.Plural är plural nu inte mer,Och söt vad bittert var innan.Vad är jag?
		-- Gopete Sherany

%
En man är som en rostig hjul på en rostig vagn,Han sjunger sin sång som han skramlar tillsammans och sedan faller han isär.
		-- Richard Thompson

%
En geni gör inga misstag.Hans fel är vilje och är portaler upptäckts.
		-- James Joyce, "Ulysses"

%
En man som fiskar efter marlin i dammarkommer att sätta sina pengar i etruskiska obligationer.
		-- James Joyce, "Ulysses"

%
En mäktig varelse är grodden,Även mindre än TJOCKHUDING.Sin vanliga bostad platsÄr djupt inne i människosläktet.Hans barnsliga stolthet han ofta behagarGenom att ge människor konstiga sjukdomar.Har du, min tallriks känner sjuka?Du innehåller förmodligen en bakterie.
		-- Ogden Nash

%
En gris är en glad följeslagare,Galt, sugga, skottkärra, eller förgylld -En gris är en kompis, som kommer att öka din moral,Även bergen kan störta och tilt.När de har blackballed, förvirrade och brände dig,När de har vänt på dig, Tory och Whig,Även om du kan kastas över av Tabby och Rover,Du kommer aldrig gå fel med en gris, en gris,Du kommer aldrig gå fel med en gris!
		-- Thomas Pynchon, "Gravity's Rainbow"

%
En robinredbreast i en burSätter alla himlen i ett raseri.
		-- Blake

%
En salamander scurries till låga för att förstöras.Imaginära varelser är fångade i födelsen på celluloid.Jag vet inte vad det handlar om. Jag är bara trummisen. Fråga Peter.föregående års Genesis utgåvan, "The Lamb Lies Downpå Broadway ".
		-- Phil Collins in 1975, when asked about the message behind

%
En enda flow'r han skickade mig, eftersom vi träffade.Alla ömt hans budbärare han valde;Djup hjärtat, ren, med doftande dagg fortfarande wet--En perfekt ros.Jag visste det språk som floweret;"Mina sköra blad", det sade, "hans hjärta bifoga."Älskar långa har tagit för hans amulettEn perfekt ros.Varför är det ingen någonsin skickade mig ännuEn perfekt limousine, tror du?Ah nej, det är alltid bara min tur att fåEn perfekt ros.
		-- Dorothy Parker, "One Perfect Rose"

%
En sanning som berättas med onda avsikterSlår alla lögner du kan uppfinna.
		-- William Blake

%
A-Z givet,1-10 alfabetiskt,härifrån till evigheten utan i betweens,fortfarande letar efter en perfekt passform i en off-the-rack världen,Försäljnings föredrag från försäljarenär allt jag vill göra är att sänka motstånd,ingen rytm i cymbaler ingen tempo i fat,kärlekens vid ankomsten,Hon kommer när hon kommer,rätt på målet, men målet i den ...
		-- William Blake

%
Abou Ben Adhem (kan hans stam öka!)Vaknade en natt från en djup dröm om fred,Och såg, i månskenet i sitt rum,Att göra det rika, och som en lilja i blom,En ängel skriver i en bok av guld.Överstiger fred hade gjort Ben Adhem fet,Och på närvaron i rummet sade han,"Vad har skrivit på du?" Visionen höjde sitt huvud,Och med en blick gjord av alla söta överenskommelseSvarade: "Namnen på dem som älskar Herren.""Och är min man?" sa Abou. "Nej inte så"Svarade ängeln. Abou talade mer låg,Men cheerly fortfarande; och sade: "Jag ber dig då,Skriv mig som en som älskar hans kolleger-män. "Ängeln skrev, och försvann. Nästa nattDet kom igen med en stor uppvaknande ljus,Och visade namnen som kärlek till Gud hade välsignat,Och lo! Ben kända Adhems ledde allt det andra.
		-- James Henry Leigh Hunt, "Abou Ben Adhem"

%
Efter ett tag lär den subtila skillnadenMellan hålla en hand och kedja en själ,Och du veta att kärlek betyder inte säkerhet,Och du börjar att lära sig att kyssar är inte kontraktOch presenterar inte löftenOch du börjar att acceptera dina förlusterMed huvudet upp och ögonen öppna,Med nåden av en kvinna, inte sorg av ett barn,Och du lär dig att bygga alla dina vägarPå dagens eftersom morgondagens jordÄr alltför oviss. Och terminer harEtt sätt för att falla ned i midflight,Efter ett tag lär att även solsken brinner om du får för mycket.Så du planterar din egen trädgård och dekorera din egen själ, i stället för att väntaFör någon att ge dig blommor.Och du lär dig att du verkligen kan uthärda ...Att du verkligen är starka,Och du verkligen har värtOch du lär och läraMed varje adjö lära dig.
		-- Veronic Shoffstall, "Comes the Dawn"

%
Efter all min dåvarande kära,Min inte längre omhuldade,Behöver vi säga att det var inte kärlek,Bara för att det dog?
		-- Edna St. Vincent Millay

%
flydde igen hon, men snabbt han kom.Tin "uviel! Tin "uviel!Han kallade henne vid hennes alviska namn;Och det stoppade hon lyssnar.Ett ögonblick stod hon, och ett passHans röst som på henne Beren komOch undergång föll på Tin "uvielAtt i sina armar låg gnistrande.Som Beren såg in i hennes ögonInom skuggorna i hennes hår,Den darrande starlight av luftrummetHan såg att det speglade skimrande.Tin "uviel Elven-mässan,Odödlig jungfru elven-wise,Om honom kastade henne skugg hårOch armar som silver glimrande.Lång var det sätt som ödet dem bar,O'er steniga berg kallt och grått,Genom hallar av järn och darkling dörr,Och skogar Nights morrowless.De Sundering Seas mellan dem låg,Och ändå till sist de möttes igen,Och länge sedan de gått bortI skogen sjunga sorrowless.
		-- J. R. R. Tolkien

%
Mot Idleness och MischiefHur förtär lite upptagen bee hur skickligt hon bygger sin cell!Förbättra varje lysande timme, hur snyggt hon sprider vaxet!Och samla honung hela dagen och mödor svårt att förvara den välFrån varje öppning blomma! Med den söta mat hon gör.I verk av arbetskraft eller skicklighet i böcker, eller arbete, eller hälsosam spel,Jag skulle vara alltför upptagen; Låt mina första år föras,För Satan finner några bus ändå att jag kan ge för varje dagFör sysslolösa händer att göra. Några bra konto till sist.
		-- Isaac Watts, 1674-1748

%
Ah, men en mans grepp bör överskrida hans räckhåll,Eller vad är ett himmelrike för?
		-- Robert Browning, "Andrea del Sarto"

%
Ah, men valet av drömmar att leva,det är där skon klämmer.För alla drömmar är inte lika,någon utgång till mardrömmest ände med drömmarenMen åtminstone en måste levas ... och dog.
		-- Robert Browning, "Andrea del Sarto"

%
Ah, mina vänner, från fängelset, frågar de till mig,"Hur bra, hur bra känns det att vara fri?"Och jag svarar dem mest mystiskt:"Är fåglar fria från kedjorna av sky-vägen?"
		-- Bob Dylan

%
Aleph-null flaskor öl på väggen,Aleph-null flaskor öl,Du tar en ner, och ge det runt,Aleph-null ölflaskor på väggen.
		-- Bob Dylan

%
Alive utan andetag,Så kallt som döden;Aldrig törstig, någonsin dricka,Sammantaget post aldrig spottar.
		-- Bob Dylan

%
Allt jag behöver ha en bra tid,Är en marijuanacigarett, en kvinna och en flaska vin.Med dessa tre saker som jag inte behöver ingen sol,En marijuanacigarett, en kvinna och en flaska vin.Allt jag vill är att aldrig bli gammal,Jag vill tvätta i ett badkar av guld.Jag vill 97 kilo redan rullat,Jag vill tvätta i ett badkar av guld.Jag vill tända mina cigarrer med 10 dollarsedlar,Jag vill ha en boskapsranch i Beverly Hills.Jag vill ha en flaska Red Eye som alltid är fylld,Jag vill ha en boskapsranch i Beverly Hills.
		-- Country Joe and the Fish, "Zachariah"

%
Alla mina vänner är gifta,Ja, de är alla bli gammal,De är alla stanna hemma på helgen,De är alla gör vad de blir tillsagda.
		-- Country Joe and the Fish, "Zachariah"

%
Allt som är guld inte glitter,Inte alla som vandrar är vilsna;Den gamla som är stark inte vissna,Djupa rötter är inte nås av frost.Ur askan en brand skall väckas,Ett ljus från skuggorna skall komma;Förnyad skall vara blad som var bruten,Den crownless igen skall vara kung.
		-- J. R. R. Tolkien

%
Allt som du trycker på, och allt du skapar,Allt som du ser, och allt du förstör,Allt som du smaka, Allt som du gör,Allt du känner, och allt du säger,Och allt som du älskar, Allt som du äter,Och allt som du hatar, och alla du möter,Allt du misstro, allt som du lätt,Allt du spara och alla du slåss,Och allt som du ger, och allt som är nu,Och allt som du behandlar, och allt som är borta,Allt som du köper, och allt som är att komma,Beg, låna eller stjäla, och allt under solen är						i samklang,Men solen förmörkasAv månen.Det finns ingen mörk sida av månen ... verkligen ... I själva verket är det allt mörkt.
		-- Pink Floyd, "Dark Side of the Moon"

%
Alla linjer har skrivits Det har varit Sandburg,Det är tråkigt, men det är sant Keats, Poe och McKuenMed alla orden borta, de hade alla deras dagVad är en ung poet att göra? Och visste vad de doin 'Men alla de ord skrivna Fågeln är en konstig en,Och alla linjer läsa, så liten och så anbudDet finns ett jag gillar mest, sin ras fortfarande okänd,Och av en fågel sades! För att inte nämna dess kön.Det påminner mig om dagar Vad är denna linjeBåde dysterhet och av ljus. Vems författarens okändDen lyfter fortfarande humöret och fortfarande gör mig fnissaOch börjar dagen på rätt sätt. Även nu när jag vuxit?Jag har läst alla de storaBåde svältande och fett,Men ingen var lika stor som"Jag tot I-taw en puddy tat."
		-- Etta Stallings, "An Ode To Childhood"

%
Hela världen är en VAX,Och alla kodare endast slaktare;De har sina utgångar och deras inälvor;Och en int i sin tid spelar många bredder,Hans sizeof väsen _ N bytes. Vid första spädbarnet,Mewling och vördnadsfull i Regent armar.Och sedan gnälla skol, med sin sol,Och lysande morgon ansikte, krypande som snigelMotvilligt till skolan.
		-- A Very Annoyed PDP-11

%
Alla som glädje skulle vinna måste dela det -Lycka föddes en tvilling.
		-- Lord Byron

%
Ett öga i en blå ansikteSåg ett öga i ett grönt ansikte."Det öga är så här öga"Sade den första ögat,"Men i låg plats,Inte i hög plats. "
		-- Lord Byron

%
En Hacker det var en av de finaste sortSom kontrollerade systemet; grafik var hans sport.En manlig man, att vara en trollkarl kan;Många en skyddad fil han sitter på sitt bord.Hans konsol, när han skrev, en man kan höraKlicka och feeping vind så tydlig,Ja, och så högt som gör maskinrummet bellDär min herre Hacker var Före av cellen.Rättsstats bra St Savage eller St DoeppnorSom gammal och strikt han tenderade att ignorera;Han släppte av de saker i gårOch tog den moderna världens rymligare sätt.Han gradera inte denna text som en plockad hönaSom säger att Hackare är inte heliga män.Och att en hacker underworked är en renFisk på torra land, flaxande på piren.Det vill säga, en hacker ut ur hans kloster.Det var en text han höll inte värt ett ostron.Och jag gick och sade hans åsikter var god;Skulle han studera till huvudet wend runtLutad över böcker i klostret? Måste han sliterSom Andy bad och ända till jorden?Skulle han lämna världen på hyllan?Låt Andy har hans arbete för sig själv![Väl, nästan. Ed.]
		-- Chaucer

%
Och allt som Lorax kvar här i den här röranvar en liten hög med stenar med ett ord, "om inte".Vad det innebar, ja, jag bara kunde inte gissa.Det var länge, länge sedan, och varje dag sedan den dagen,Jag har orolig och bekymrad och orolig bort.Genom åren som mina byggnader har fallit isär,Jag har orolig det med hela mitt hjärta."Men", säger Oncler, "nu när du är här,ord Lorax verkar helt klart!Om inte någon som du bryr sig hela massa,ingenting kommer att bli bättre - det är inte.Så ... fångst! "Ropar Oncler. Han låter något fall."Det är en Truffula frö. Det är den sista av alla!"Du är ansvarig för den sista av de Truffula frön.Och Truffula träd är vad alla behöver.Plantera ett nytt Truffula - behandla den med omsorg.Ge det rent vatten och mata den friska luften.Odla en skog - skydda den från axlar som hacka.Då Lorax och alla hans vänner kan komma tillbaka! "
		-- Chaucer

%
Och som vi står på kanten av mörkerLåt vår sång fylla tomrummetAtt andra kan kännaI landet i nattenFartyget av solenDras avDen tacksamma döda.
		-- Tibetan "Book of the Dead," ca. 4000 BC.

%
Och gjorde dessa fötter, i gamla tider,Gå på Englands berg grönt?Och var den Helige Guds LammI Englands trevliga betesmarker sett?Och gjorde Skepnaden gudomligaLysa på dessa trångt kullar?Och var Jerusalem byggde härBland dessa mörka sataniska fabriker?Ge mig min båge av brinnande guld!Ge mig mina pilar av lust!Ge mig mina spjut! O moln utvecklas!Ge mig min vagn av eld!Jag ska inte upphöra av psykisk kamp,Inte heller skall mitt svärd vila i min hand,Tills vi har byggt JerusalemI England gröna och angenäma land.
		-- William Blake, "Jerusalem"

%
Och här jag vänta så tålmodigtVäntar på att ta reda på vad prisDu måste betala för att få ut avGår igenom alla dessa saker två gånger
		-- Dylan, "Memphis Blues Again"

%
Och jag hörde Jeff utbrista,När de vandrade ut ur sikte,"God jul till alla -Du tar kreditkort, eller hur? "
		-- "Outsiders" comic

%
Och om Kalifornien glider ut i havet,Liksom mystiker och statistik säger att det kommer.Jag förutspår denna Motell kommer att stå,Tills jag har betalat min räkning.
		-- Warren Zevon, "Desperados Under the Eaves"

%
Och om någon gång, någonstans, beder någon dig,"Vem kilt dig?", Berätta det Twas Doones av Bagworthy!
		-- Warren Zevon, "Desperados Under the Eaves"

%
Och om du undrar,Vad jag gör,Som jag är på väg för sink.Jag spottar ut all bitterhet,Tillsammans med hälften av min sista drink.
		-- Warren Zevon, "Desperados Under the Eaves"

%
Och i Heartbreak år som ligger framför oss,Var sann mot dig själv och Grateful Dead.
		-- Joan Baez

%
Och miles för att gå innan jag sover.
		-- Robert Frost

%
Och nu din toner är toney, Disk block aplentyOch papperet nära ren vit, väntar på ditt laser dras linjer,De fläckar på din själ är borta Dina intrikata typsnitt,Och utskrifterna är ren så lätt .. Dina bilder och tecken.Vi har arbetat med din far, din amputative frånvaroDen ärevördiga XGP, har gjort tio dum,Men hans långsamma konstnärliga handen, Utan dig, Dover,Saknar din ren hastighet. Vi är systemet untounged-Avhandlingar och uppsatser DRAW täppor och TEXageOch kod i en kö Har bidade sin tid,Dover, oh Dover, med LISP kod och program,Vi har väntat på dig. Och detta crufty rim.Dover, oh Dover, Dover, oh Dover, uppstått från döda.Vi välkomnar dig tillbaka, Dover, oh Dover, vaknat ur sängen.Men fortfarande kan du fastna, Dover, oh Dover, välkommen tillbaka till labbet.Du är på rätt spår. Dover, oh Dover, har vi missat din renahand ...
		-- Robert Frost

%
... och rapportkort Jag var alltid rädd för att visaMama'd komma till skolanoch som jag skulle sitta där mjukt CryinTeacher'd säger att han är bara inte tryin 'Fick ett bra huvud om han skulle tillämpa detmen du känner dig självDet är alltid någon annanstansJag skulle bygga mig ett slottmed drakar och kungaroch jag skulle åka ut med demNär jag stod vid mitt fönsteroch såg ut på deBrooklyn vägar
		-- Neil Diamond, "Brooklyn Roads"

%
Och så var det senare,Som mjölnaren berättade sin historia,Att hennes ansikte, först bara spöklikt,Vände en vitare nyans av blek.
		-- Procol Harum

%
Och tystnaden kom böljande mjukt bakåtNär störtar hovar var borta ...
		-- Walter de La Mare, "The Listeners"

%
Och det är bra gamla Boston,Hemma hos bönor och torsk,Där Lowells tala endast Cabots,Och Cabots prata bara till Gud.
		-- Walter de La Mare, "The Listeners"

%
Och vi hörde honom utropaNär han började ströva:"Jag är ett hologram, barn,försök inte detta hemma! "
		-- Bob Violence

%
Och ... Vad händer i världen någonsin blev Sweet Jane?Hon har förlorat sin gnistan, ser att hon är inte samma sak.Livin på reds, C-vitamin, och kokainAllt en vän kan säga är "Är det inte synd?"
		-- The Grateful Dead

%
Änglar vi har hört på högBerätta att gå ut och köpa.
		-- Tom Lehrer

%
Antonio AntonioVar trötta på att leva alonioHan trodde att han skulle uppvakta Antonio AntonioMiss Lucamy Lu, Rode av hans polo ponioMiss Lucamy Lucy Molonio. Och hittade piganI en bowery skugga,Sitter och stickning alonio.Antonio AntonioSagt om du blir min ownioJag kommer att älska tou sant Oh Nónio AntonioOch köp för dig Du är alldeles för dyster och bonioEn icery creamry Conio. Och allt som jag önskarDu singular fiskÄr att du snabbt kommer begonio.Antonio AntonioYttrade en dyster moanioOch gick och gömdeEller jag höra att han gjordeI Antartical Zonio.
		-- Tom Lehrer

%
April är den grymmaste månaden ...
		-- Thomas Stearns Eliot

%
Finns det sådana i landet av de modigaVem kan berätta för mig hur jag ska beteNär jag vanäradeEftersom jag raderadeEn fil jag tänkt att spara?
		-- Thomas Stearns Eliot

%
När det gäller kvinnor, men vi hånar och struntar dem,Vi kan leva med, men kan inte leva utan dem.
		-- Frederic Reynolds

%
Som jag gick upp hålkort Hill,Känsla värre och värre,Där träffade jag en C.R.T.Och det drop't mig en markör.C.R.T., C.R.T.,Fosfor ljus på dig!Om jag hade femtio timmar per dagJag skulle spendera dem alla på dig.
		-- Uncle Colonel's Cursory Rhymes

%
Som jag passerar Project MAC,Jag träffade en Quux med sju hacka.Varje hacka hade sju buggar;Varje bugg hade sju manifestationer;Varje manifestation hade sju symptom.Symptom, manifestationer, buggar, och hackar,Hur många förluster på Project MAC?
		-- Uncle Colonel's Cursory Rhymes

%
Som jag gick ner på gatan en mörk och trist dag,Jag kom på en skylt och mycket till min bestörtning,Orden var rivna och sliten,Från stormen natten innan,Vind och regn hade gjort sitt arbete och detta är hur det går,Rök Coca-Cola cigaretter, tugga Wrigleys Spearmint öl,Ken-L-Ration hundmat gör din hy klar,Simonize ditt barn i en Hershey candy bar,Och Texaco är en skönhet grädde som används av varje stjärna.Ta din nästa semester i en helt ny Frigedaire,Lära sig att spela piano i vinter underkläder,Läkare säger att barn ska röka tills de är tre,Och personer över sextiofem bör bada i Lipton te.
		-- Uncle Colonel's Cursory Rhymes

%
Som mig en "mig marrer var Readin en tyape,Den tyape gav ett skrik markera ett "försökt tae escyape;Det hoppas över ower den gyate tae slutet av fältet,En "pimplas oot rummet wi" en spole en "en rulle!Följ ledare, Johnny mig laddie,Följer den genom, me slug lad O;Följ transport, Johnny mig laddie,Bort, gosse, ligger bort, slug lad O!
		-- S. Kelly-Bootle, "The Devil's DP Dictionary"

%
Som en dag kan det hända att ett offer måste hittasJag har en liten lista - Jag har en liten listaSamhällets brottslingar som kan mycket väl vara under jordOch som aldrig skulle missas - som aldrig skulle missas.
		-- Koko, "The Mikado"

%
Ibland diskretion bör kastas åt sidan,och med den dåraktiga ska vi spela idiot.
		-- Menander

%
Undvik Tyst och Placid personer om du inte är i behov av sömn.
		-- National Lampoon, "Deteriorata"

%
Azh nazg durbatal ^ uk, azh nazg gimbatul,Azh nazg thrakatal ^ uk agh burzum ishi krimpatul!
		-- J. R. R. Tolkien

%
Vara säker på att en promenad genom havet av de flesta Souls skulle knappastfå dina fötter är våta. Fall inte in Love, därför: det kommer att hålla i ansiktet.
		-- National Lampoon, "Deteriorata"

%
Vara tapper, men inte alltför VÅGHALSIG.Låt din klädsel vara comely, men inte kostsamt.
		-- John Lyly

%
Skönhet är sanning, sanning skönhet, det är alltVeten på jorden, och alla ni behöver veta.
		-- John Keats

%
Eftersom jag gör,Eftersom jag inte hoppas,Eftersom jag inte hoppas att överlevaOrätt från slottet, död från luften,Eftersom jag bara göra,Jag fortsätter...
		-- T. S. Pynchon

%
Under denna sten ligger Murphy,De begravde honom i dag,Han levde livet av Riley,Medan Riley var borta.
		-- T. S. Pynchon

%
rop bättre! lyra!bättre watchoutlpr varförjultomten <nordpolen> stadcat / etc / passwd> listannKontrollera listanKontrollera listacat lista | grep stygg> nogiftlistcat lista | grep trevligt> Gåvolistajultomten <nordpolen> stadsom | grep sovandesom | grep vakensom | grep "dåliga \ | bra"	för Guds skull) {		var snäll}
		-- T. S. Pynchon

%
Mellan idénOch verklighetenMellan rörelseOch lagenFaller Shadow[Citerat i "VMS interna och datastrukturer", V4.4, närmed hänvisning till systemtjänstexport.]
		-- T. S. Eliot, "The Hollow Man"

%
Big M, Little M, många mumlande mössGör midnatt musik i månskenet,Mighty nice!
		-- T. S. Eliot, "The Hollow Man"

%
Bit utanför mer än mitt sinne kunde tugga,Dusch eller självmord, vad ska jag göra?
		-- Julie Brown, "Will I Make it Through the Eighties?"

%
Svart glänsande Molly och ljusa färgade guppy,Shy små änglar så skonsam som valpar,Simning och dykning med knappt en sus,De var bara några av mina tropiska fiskar.Sen fick jag mantor som sticker i vattnet,Dödliga pirayor som kliar för en slakt,Savage manliga beta som biter med en squish,Nu har jag många mindre tropiska fiskar.Om du tror attFisk är fredligaDet är ett tomt önskan.Bara dumpa dem tillsammansOch lämna dem ifred,Och snart kommer du att ha - ingen fisk.
		-- To My Favorite Things

%
Blackout, värmebölja, 0,44 kaliber mord,Bums drop dead och hundarna galen i förpackningar på västra sidan,En ung flicka som står på en avsats, ser ut som en annan självmord,Hon vill träffa dessa tegelstenar,"Orsaka att nyheterna på sex fick hålla sig till en deadline,Medan miljonärer gömma sig i Beekman plats,De väska damer kastar sina ben i ansiktet,Jag blir attackerad av en unge med stereoljud,Jag vill inte höra det, men han kommer inte att stänga ner ...
		-- Billy Joel, "Glass Houses"

%
Pojke, få huvudet ur stjärnorna ovan,Du får maximal glädje av ett minimum av kärlek.Spara ditt hjärta och låta kroppen vara tillräckligt,För att få maximal glädje av ett minimum av kärlek.Spara ditt hjärta och låta kroppen vara tillräckligt,Och få maximal glädje av ett minimum av kärlek.
		-- Mac Macinelli, "Minimum Love"

%
Andas djupt insamling dysterhet.Titta ljus bleknar från varje rum.Säng-sitter människor ser tillbaka och klagan;en annan dagens värdelös energier spenderas.Passionerade älskande brottas som en.Ensam man ropar efter kärlek och har ingen.Ny mamma plockar upp och diar sin son.Pensionärer önskar att de var unga.Kallsinnig orb som härskar natten;Tar bort färger från vår syn.Rött är grå och gul vit.Men vi avgöra vilka är verkliga, och som är en illusion. "
		-- The Moody Blues, "Days of Future Passed"

%
Brillineggiava, ed i tovoli slatigirlavano ghimbanti nella vaba;Jag borogovi eran tutti mimantie la moma radeva fuorigraba."Figliuolo mio, sta" Attento al Gibrovacco,dagli artigli e dal Morso lacerante;Fuggi l'uccello Giuggiolo, e nel SaccoMetti infine il frumioso Bandifante ".
		-- Lewis Carroll, "Jabberwocky"

%
Men har någon liten atom,Medan a-sittin 'och en-splittin',Någonsin slutat tänka eller CAREAtt E = m c ** 2?
		-- Lewis Carroll, "Jabberwocky"

%
Men jag var där och jag såg vad du gjorde,Jag såg det med mina egna två ögon.Så du kan torka bort det grin;Jag vet var du har been--Det är allt varit en lögn!
		-- Lewis Carroll, "Jabberwocky"

%
Men forskarna, som borde vetaFörsäkra oss om att det måste vara så.Åh, låt oss aldrig, aldrig tvivelVad ingen är säker på.
		-- Hilaire Belloc

%
Men mjuk du det verkliga Ophelia:Ope icke dina otympliga och marmor käftar,Men få dig till ett nunnekloster - gå!
		-- Mark "The Bard" Twain

%
Men, Mousie, du är ingen din körfält,Bevisa förutseende kan vara förgäves:De bästa som system o 'möss en "mänGang akter a-gley,En "lea'e oss intet annat än sorg och smärtaFör utlovade glädje.
		-- Robert Burns, "To a Mouse", 1785

%
Surrar av, banan näsa; Lindra mina ögonAv hatiskt ömhet, rensa mina ax;Mindre kär än armémyror i äppelpajerDu, gamla beskära ansikte, med dina kastanjer slitna,Dropt från din peeling läppar som usel frukt;Liknande honungsbin på de överlämnade perfum'd ökadeDe suger och gillar dubbelknäppt kostymÄr inaktuell; Därför, banan näsa,Gå flyga drake, din välkomna är overstayed;Och hejda produkter av dina waspish förstånd:Thy logick, likt ditt lås, är disarrayed;Din jubel, liksom din hy, är gropar.Var off säger jag; gå bugg någon ny,Snabbstopp, slå det, få dig därmed och nötter till dig.
		-- Robert Burns, "To a Mouse", 1785

%
Vid tiden du svär du är hans,frossa och suckandeoch han lovar hans passion äroändlig, odödliga -Lady, anteckna detta:En av er ligger.
		-- Dorothy Parker, "Unfortunate Coincidence"

%
Genom gården, livet är hårt.Genom tum, är det en enkel match.
		-- Dorothy Parker, "Unfortunate Coincidence"

%
Lugna ner, det är bara ettor och nollor,Lugna ner, det är bara bits och bytes,Lugna ner och prata med mig på engelska,Vänligen inse att jag inte är en av dina computerites.
		-- Dorothy Parker, "Unfortunate Coincidence"

%
Avbryt mig inte - för vad då skall förbli?Abskissan vissa mantissorna, moduler, lägen,En rot eller två, en torus och en nod:Inversen av min vers, en noll domän.
		-- Stanislaw Lem, "Cyberiad"

%
Godisär dandymen spritÄr snabbare.Fortune uppdaterar stora citat: # 53.Candy är dandy; men sprit är snabbare,och kön inte kommer att ruttna tänderna.
		-- Ogden Nash, "Reflections on Ice-Breaking"

%
Fånga en våg och du sitter på toppen av världen.
		-- The Beach Boys

%
Cecil, du är mitt sista hoppAtt ta reda på den verkliga Straight DopeFör jag har läst av Schrödingers kattMen ingen av mina katter inte alls så.Denna ovanliga djur (så sägs det)Är samtidigt levande och död!Vad jag inte förstår är varför just hanKan inte vara det ena eller det andra, utan tvekan.Min framtid hänger nu mellan egentillstånd.I en Jag är upplyst, i det andra jag inte.Om * du * förstå, Cecil, visa mig då vägenOch rädda mitt psyke från kvant förfall.Men om queer sak har förbryllat även du,Då ska jag * ___ och * Jag kommer inte att se dig i Schrodingers zoo.av mänsklig kunskap "av Cecil Adams
		-- Randy F., Chicago, "The Straight Dope, a compendium

%
Visst finns det saker i livet som pengar kan inte köpa,Men det är väldigt roligt - har du någonsin försöka köpa dem utan pengar?
		-- Ogden Nash

%
Charlie var en kemist,Men Charlie är inte mer.För vad han trodde var H2O,Var H2SO4.
		-- Ogden Nash

%
Barn är inte nöjda utan något att ignorera,Och det är vad föräldrarna skapades för.
		-- Ogden Nash

%
Ridderlighet, Schmivalry!Roger tjuven har enmetod han använder förlömsk attacker:Folk som läser ärkarakteristisktAlltid glömmer attVakta sin egen bac ...
		-- Ogden Nash

%
Jultid är här, vid Golly; Döda kalkoner, ankor och höns;Ogillande skulle vara dårskap; Blanda stansen, dra ut Dickens;Deck the halls med hunks av järnek, Även om utsikterna sickens,Fyll koppen och inte säga när ... Brother, här går vi igen.På juldagen, kan du inte få ont; Förbindelser spara några expense'll,Din medmänniska måste du älskar; Skicka några värdelös gamla redskap,Det är dags att råna honom allt mer, eller en matchande penna och penna,De övriga 364! Bara det jag behöver ... hur trevligt.Det spelar ingen roll hur uppriktig Hark The Herald-Tribune sjunger,Det är inte heller hur innerlig anden; Reklam fantastiska saker.Känslan kommer inte att göra kär den; God Rest Ye Merry Merchants,Vad som är viktigt är ... priset. Kan du göra Yuletide lön.Änglar som vi har hört på High,Låt vild Sleigh Bells jingle; Berätta att gå ut och köpa.Hagel vår kära gamla vän, Kris Kringle, Sooooo ...Kör sin renar över himlen,Stå inte under när de flyger förbi!
		-- Tom Lehrer

%
Kall för hand och hjärta och ben,och kall vara sova under sten;aldrig mer att vakna på stenig säng,aldrig, tills solen misslyckas och månen är död.I den svarta vinden stjärnorna skall dö,och fortfarande på guld här låta dem ligga,till den mörka herre lyfter sin handöver döda havet och vissnade land.
		-- J. R. R. Tolkien

%
Kom och fyll koppen och eld vårenDin vinterplagg av ånger fling.Fågeln tid har men en liten vägFladdra - och fågeln är på vingen.
		-- Omar Khayyam

%
Bo hos mig och vara min kärlek,Och vi kommer vissa nya nöjen bevisaAv gyllene sand och kristall bäckarMed silkes linjer och silver krokar.Det finns ingenting som jag inte skulle göraOm du vill bli min POSSLQ.Du bor med mig, och jag med dig,Och du kommer att bli min POSSLQ.Jag vill vara din vän och så mycket mer;Det är vad en POSSLQ är för.Och allt kommer vi att erkänna;Ja, till och med IRS.En dag på vad vi båda kan tjäna,Kanske kommer vi att lämna in en gemensam avkastning.Du kommer att dela min pad, min skatt, joint;Du kommer att dela mitt liv - upp till en punkt!Och att du kommer att bli så glad att göra,Eftersom du kommer att bli min POSSLQ.
		-- Omar Khayyam

%
Bo hos mig, och vara min kärlek,Och vi kommer vissa nya nöjen bevisaAv gyllene sand och kristall bäckar,Med silkes linjer och silver krokar.
		-- John Donne

%
Kom igen, Virginia, gör inte mig vänta!Katolik flickor börjar alldeles för sent,Ah, men förr eller senare kommer det ner till ödet,Jag kan lika gärna vara en.Tja, visade de en staty, sagt att be,Byggt ett tempel och låst bort dig,Ah, men de har aldrig sagt det pris som du har betalat,De saker som du kan ha gjort.Så kom igen, Virginia, visa mig ett tecken,Skicka upp en signal, jag ska kasta dig en linje,Som målat glas gardin som du gömmer sig bakom,Aldrig släpper in solen.Darling, bara bra dör unga!
		-- Billy Joel, "Only The Good Die Young"

%
Kom, längtar varje stympad att vara en kon,Och varje vektor drömmar om matriser.Hör till den milda lutning vinden:Det viskar av en mer ergodisk zon.
		-- Stanislaw Lem, "Cyberiad"

%
Kom, hyresvärd, fylla den strömmande skål tills det löper över,Ikväll kommer vi alla glatt vara - i morgon kommer vi att få nykter.
		-- John Fletcher, "The Bloody Brother", II, 2

%
Kom, låt oss skynda till ett högre plan,Där dyader trampa fairy områdena Venn,Sina index bedecked från en till _ n,Blandas i en ändlös Markov kedja!
		-- Stanislaw Lem, "Cyberiad"

%
Kom, musa, låt oss sjunga om råttor!
		-- From a poem by James Grainger, 1721-1767

%
Kom, ni spritSom tenderar på dödliga tankar, Unsex mig här,Och fylla mig, från kronan till tå, topp fullAv direst grymhet! göra tjock mitt blod,Stoppa upp tillgången och passagen till ångerAtt ingen compunctious besöker naturSkaka min föll ändamål, inte hålla fred mellanEffekten och det! Kom till min kvinnans bröst,Och ta min mjölk för galla, du mörda ministrar,Oavsett var i din blinda ämnenDu väntar på naturens bus! Kom, tjock natt,Och Pall den i dunnest röken av helvetet,Att min skarp kniv ser inte såret det gör,Nor himmel kika genom täcket av den mörka,Att gråta `Håll, håll!
		-- Lady MacBeth

%
Kommer till butiker nära dig:101 Grammatically Rätt Populära Tunes Presentera:(Du är inte något annat än en) Hound DogDet betyder inte en sak om det inte har fått Det SwingJag inte FelaktigtOch en hel del mer ...
		-- Lady MacBeth

%
Förvirring kommer att bli min epitafiumnär jag går en sprucken och bruten banaOm vi ​​gör det kan vi alla sitta tillbaka och skrattamen jag är rädd att vi i morgon kommer att gråta.
		-- King Crimson, "In the Court of the Crimson King"

%
Döden kommer på varje passerande vind,Han lurar i varje blomma;Varje årstid har sin egen sjukdom,Dess fara - varje timme.
		-- Reginald Heber

%
Däck oss alla med Boston Charlie,Walla Walla, Washington., En "Kalamazoo!Noras Freezin på vagnen,Swaller dollar blomkål, alleygaroo!Gör vi inte vet föråldrade fat,Vaggvisa Lilla pojke, Louisville Lou.Trolley Molly inte älskar Harold,Boola Boola Pensacoola hullabaloo!
		-- Pogo, "Deck Us All With Boston Charlie" [Walt Kelly]

%
Förklaras skyldig ... att visa känslor av en nästan mänskliga naturen.
		-- Pink Floyd, "The Wall"

%
Despising maskiner till en människa,Den Luddites gick med Klanen,Och rida ut på nattenI ett arkmaterial enligt vitLynch alla robotar de kan.
		-- C. M. and G. A. Maxson

%
Didja "någonsin måste göra upp dig,Plocka upp en och lämna andra bakom,Det är inte ofta lätt, och det är inte ofta slag,Didja "någonsin att bestämma dig?
		-- Lovin' Spoonful

%
Desillusionerade ord som kulor bark,Som mänskliga gudar sikta på sitt varumärke,Gör allt från leksakspistoler som gnistaTill hudfärgade kristusar som lyser i mörkret.Det är lätt att se utan att titta för långtAtt inte mycket är riktigt heligt.
		-- Bob Dylan

%
Gör dina utter göra shimmy?Har de gillar att skaka sina svansar?Gör dina Wombats sova i tophats?Är din trädgård full av sniglar?
		-- Bob Dylan

%
Var inte orolig, det kommer inte att skada dig,Det är bara jag fullfölja något jag är inte säker på,Över mina drömmar, med neptive konstigt,Jag jagar den ljusa svårfångade fjärilen av kärlek.
		-- Bob Dylan

%
Låt inte ingen berätta vad du inte kan göra;låt inte ingen berätta vad som är omöjligt för dig;låt inte ingen berätta vad du måste göra,eller att du aldrig vet ... vad som finns på andra sidan av regnbågen ...kom ihåg, om du inte följer dina drömmar,du vet aldrig vad som finns på andra sidan av regnbågen ...
		-- melba moore, "the other side of the rainbow"

%
Tappa inteDitt huvudFör att få en minutDu behöver ditt huvudDin hjärna är i det.
		-- Burma Shave

%
Inte väcka mig upp för tidigt ...Ska ta en tur över månen ...Du och jag.
		-- Burma Shave

%
Dubbel Bucky, du är en,Du gör mitt tangentbord så mycket kul,Dubbel Bucky, en extra bit eller två, (Vo-vo-de-o)Kontroll och meta, sida vid sida,Augmented ASCII, 9 bitar bred!Dubbel Bucky, en halv tusen tecken, plus några!Åh, jag säker önskar att jag,Hade ett par bitar mer!Kanske en uppsättning pedaler för att göra antalet bitar fyra.Dubbel Bucky! Dubbel Bucky vänster och högerOR'd tillsammans, outta syn!Dubbel Bucky, jag vill ha en hel ord,Dubbel Bucky, jag är glad att jag hört talas om,Dubbel Bucky, jag vill ha en helt ord av dig!läggas till terminalkoder på 36-bitars maskiner för användningav skärm redaktörer. [Till tonerna av "Rubber Ducky"]
		-- to Nicholas Wirth, who suggested that an extra bit

%
Ner till bananrepubliker,Ner till tropisk sol.Gå de bosatta utomlands amerikaner,I hopp om att hitta lite kul.Några av dem gå för segling,Fångas av drag av havet.Försöker hitta vad som är sjuklig,Bor i landet av den fria.Några av dem kör från vänner,Lämnar inga framåtadress.Några av dem kör massor av ganja,Vissa kör från IRS.Sent på kvällen hittar dem,I billiga hotell och barer.Stressade de senoritas,Medan de dansar under stjärnorna.
		-- Jimmy Buffet, "Banana Republics"

%
Dricka och dansa och skratta och lögnKärlek, upprullnings midnatt genomFör i morgon ska vi dö!(Men, tyvärr, vi aldrig göra.)
		-- Dorothy Parker, "The Flaw in Paganism"

%
Lätt att komma och lätt går,vissa kallar mig lätta pengar,Ibland är livet är fullt av skratt,och ibland är det inte roligtDu kanske tror att jag är en idiotoch ibland det är sant,Men jag goin 'till himlen i en blixt av brand,	med eller utan dig.
		-- Hoyt Axton

%
Eleanor RigbySitter vid tangentbordetOch väntar på en linje på skärmenBor i en drömVäntar på en signalAtt hitta någon kodDet kommer att göra maskinen göra lite mer.Vad är det för?Alla ensamma användare, var kommer de alla ifrån?Alla ensamma användare, varför tar det så lång tid?hacker MackensieSkriva koden för ett program som ingen kommer att köraDet är nästan klarTitta på honom arbeta, om fastställande av buggar i natten när det finnsingen där.Vad bryr han sig?Alla ensamma användare, var kommer de alla ifrån?Alla ensamma användare, varför tar det så lång tid?Ah, titta på alla ensamma användare.Ah, titta på alla ensamma användare.
		-- Hoyt Axton

%
Endless världens tur, oändliga solens spinningOändliga strävan;Jag vänder igen, tillbaka till min egen början,Och här, finna vila.
		-- Hoyt Axton

%
Es Brilig krig. Die Schlichte TovenWirrten und wimmelten i Waben;Und aller-m "umsige BurggovenDir mohmen R "ath ausgraben.
		-- Lewis Carrol, "Through the Looking Glass"

%
Euch ist bekannt, var wir beduerfen;Wir wollen skarp Getraenke schluerfen.
		-- Goethe, "Faust"

%
Även en man som är ren i hjärtat,Och säger att hans böner på nattenKan bli en varg när wolfbane blommar,Och månen är full och ljus.
		-- The Wolf Man, 1941

%
Även i ögonblicket då vår tidigaste kyss,När suckade ansträngt knopp i blomman,Satt torr säd mest ovälkommen detta;Och att jag visste, men inte den dagen och timmen.Alltför säsong Mässigt är jag, som land-uppfödda,Att luta på hösten eller trotsar frost:Snusning kylan även som mina fäder,Jag säger med dem, "Vad är i kväll är förlorad."Jag bara hoppades, med den milda hopp om allaSom tittar bladet ta form på trädet,En rättvisare sommaren och en senare nedgångÄn i dessa delar en man är benägen att se,Och soliga kluster mogna för vin:Jag säger er över blackened vinstockar.Vår Tidigast Kiss ", 1931
		-- Edna St. Vincent Millay, "Even in the Moment of

%
Någonsin Onward! Någonsin Onward!Det är sprit som har fört oss fame.Vi är stora men större vi blir,Vi kan inte misslyckas för alla kan se, att för att tjäna mänsklighetenHar varit vårt mål.Våra produkter nu kända i varje zon.Vårt rykte gnistrar som en pärla.Vi har kämpat oss igenomOch nya områden vi är säkra på att erövra ocksåFör någonsin Onward IBM!
		-- Ever Onward, from the 1940 IBM Songbook

%
Ända sedan jag var en ung pojke,Jag har hackat ARPA nätet,Från Berkeley ner till Rutgers, är han på min favorit terminal,Någon tillgång jag kunde få, Han katter C rakt in foo,Men inte sett något liknande honom, hans lärjungar leda honom,På varje campus ännu, och han bara bryter roten,Det döva, stumma och blinda barn, har alltid fullt SYS-PRIV-talet,Säker skickar en genomsnittlig paket. Aldrig använder ludd,Det döva, stumma och blinda barn,Säker skickar en genomsnittlig paket.Han är en UNIX-guidenDet måste finnas en snodd.UNIX guiden har är inte fick några distraktioner,Obegränsat utrymme på disken. Kan inte höra några visselpipor eller klockor,Hur tror du att han gör det? Det går inte att se något meddelande blinkar,jag vet inte. Typer av luktsinne,Vad gör honom så bra? Dessa galna små program,De korrekta bit flaggor inställd,Det döva, stumma och blinda barn,Säker skickar en genomsnittlig paket.
		-- UNIX Wizard

%
Varje kärlek är kärlek innanI en mattare klänning.
		-- Dorothy Parker, "Summary"

%
Varje människa är som Gud gjorde honom, ay, och ofta värre.
		-- Miguel de Cervantes

%
Varje natt mina böner jag säger,Och få min middag varje dag;Och varje dag som jag har varit bra,Jag får en orange efter mat.Barnet som inte är rent och snyggt,Med massor av leksaker och saker att äta,Han är en stygg barn, jag är sure--Annars hans kära pappa är dålig.
		-- Robert Louis Stevenson

%
Alla vet att tärningen är laddade. Alla rullar med derashåll tummarna. Alla vet kriget är över. Alla vet attgoda förlorade. Alla vet kampen fastställdes: den dåliga vistelsenfattiga, de rika blir rika. Det är hur det går. Alla vet.Alla vet att båten läcker. Alla vet kaptenenlied. Alla fick denna brutna känsla som sin far eller sin hundjust dött.Alla pratar med sina fickor. Alla vill ha en chokladaskoch lång stjälk ros. Alla vet.Alla vet att du älskar mig, baby. Alla vet att du verkligendo. Alla vet att du har varit trogen, ge eller ta en natt ellertvå. Alla vet att du har varit diskret, men det fanns så många människordu bara hade att möta utan dina kläder. Och alla vet.Och alla vet att det är nu eller aldrig. Alla vet att det är jag eller du.Och alla vet att du leva för evigt när du har gjort en rad eller två.Alla vet affären är ruttet: Old Black Joe fortfarande Pickin bomullför dig band och rosetter. Och alla vet.
		-- Leonard Cohen, "Everybody Knows"

%
Allt är stor i denna gamla goda världen;(Detta är saker som de kan alltid använda.)Guds i sin himmel, kullens dagg pärlgryn;(Detta kommer att ge barnets skor.)Hunger och krig betyder inte ett ting;Allt är rosen where'er vi strövar;Hark, hur småfåglarna glatt sjunga!(Detta är vad hämtar bacon hem.)
		-- Dorothy Parker, "The Far Sighted Muse"

%
Vart du än går ser du dem att söka,Överallt kommer du att känna smärta,Alla är ute efter svaret,Väl titta igen.
		-- Moody Blues, "Lost in a Lost World"

%
F: När i ett rum som jag störta, jagIbland hittar några VIOLETT svampar.Då jag kvar, mörkt grubbelPå giftet de är vätskande.
		-- The Roguelet's ABC

%
Familjer, när ett barn födsVill att det ska vara intelligent.Jag, genom intelligens,Efter att ha havererade hela mitt liv,Bara hoppas att barnet kommer att visaOkunniga och dumma.Då kommer han kröna en lugn livGenom att bli en minister
		-- Su Tung-p'o

%
Farväl vi kallar till härden och hall!Även vind kan blåsa och regnet kan falla,Vi måste bort ere rast på dagenLångt över trä och berg hög.Till Vattnadal, där alver ännu uppehållaI gläntor under dimmiga föll,Genom hed och avfall rider vi i all hast,Och vart kan vi inte tala om.Med fiender framåt, bakom oss fruktar,Under himlen ska vara vår säng,Till sist vår slit föras,Vår resa gjort, rusade vår ärende.Vi måste bort! Vi måste bort!Vi rider före paus på dagen!
		-- J. R. R. Tolkien

%
Felix Catus är din taxonomiska nomenklatur,En endotermisk quadroped, köttätande av naturen.Dina visuella, lukt- och hörsel sinnenBidra till din jakt färdigheter och naturliga försvar.Jag befinner mig fascinerad av din sub-sång svängningar,En sällsam utveckling av kattkommunikationSom undanröjer din grundläggande hedonistiska predelectionFör en rytmisk stryker av pälsen för att visa tillgivenhet.En svans är helt avgörande för dina akrobatiska talanger:Du skulle inte vara så smidig om du saknade sin motvikt;Och när den inte utilitized för att underlätta förflyttning,Det tjänar ofta för att illustrera läget i dina känslor.Oh Ställe, komplexa nivåer av beteende som du visarBeteckna en ganska väl utvecklad kognitiv array.Och om du inte är kännande, Spot, och inte förstå,Jag ändå anser dig en sann och uppskattad vän.
		-- Lt. Cmdr. Data, "An Ode to Spot"

%
Femton män på en död mans kista,Yo-ho-ho och en flaska med rom!Flaskan och fan hade gjort för resten,Yo-ho-ho och en flaska med rom!
		-- Stevenson, "Treasure Island"

%
Femtio lättvindiga grodorPromenerade genom på flippered fötterOch med sin slem de gjorde tidOnaturligt flotta.
		-- Stevenson, "Treasure Island"

%
Slutgiltig är döden.Perfektion är slutgiltig.Ingenting är perfekt.Det finns klumpar i den.
		-- Stevenson, "Treasure Island"

%
Fem namn som jag kan knappt stå att höra,Inklusive ditt och mitt och ett mer schimpansen som inte är här,Jag kan se damerna prata hur tiderna är Getting hårt,Och det skräckinjagande utgrävning på Magnolia boulevard,Ja, jag goin 'galen,Och jag skrattar åt den frusna regn,Tja, jag är så ensam, honung när de ska skicka hem mig?Dåliga gymnastikskor och en pina colada min vän,Stoppa på Avenyn med Radio City, med enTransistor och en stor summa pengar att spendera ...Du fellah, du Tearin "upp på gatan,Du bär den vita smoking, hur ska du slå värmen,Tar du mig för en idiot, tror du att jag inte ser,Det dike i dalen att de är Diggin bara för mig,Ja, och det som händer galen,Du vet att jag laughin "på den frusna regn,Känns som jag är så ensam, honung när de ska skicka hem mig?(kör)
		-- Bad Sneakers, "Steely Dan"

%
Flygande tefat på gångVisa sig att det mänskliga ögat.Aliens rök, skjuta upp invasionenMedan de profilera dessa berättelser som lögner.
		-- Bad Sneakers, "Steely Dan"

%
"För ett par O stift", säger Troll och grinar,"Jag ska äta dig också, och gnaga dina smalbenen.En bit o 'färskt kött kommer att gå ner söt!Jag ska försöka mina tänder på dig nu.Hee nu! Se nu!Jag är trött o gnagande gamla ben och skinn;Jag har lust att äta på dig nu. "Men precis som han trodde att hans middag fångades,Han fann händerna hade tag i intet.Innan han kunde tänka, Tom gled behingOch gav honom skon Lärn honom.	Varna honom! Darn honom!En bula o 'the boot på sätet, thoguht Tom,Skulle vara ett sätt att Lärn honom.Men hårdare än sten är kött och benAv ett troll som sitter i ensam kullar.Samt ställa in start till berget rot,För säte ett troll inte känna det.Skal det! Läka det!Old Troll skrattade, när han hörde Tom stöna,Och han visste att hans tår kunde känna det.Tom ben är spel, eftersom hemmet han kom,Och hans mufflös fot är bestående lama;Men Troll bryr sig inte, och han är fortfarande kvarMed benet han urbenat från sin ägare.Doner! Tabbe!Troll gamla säte är fortfarande densamma,Och benet han urbenat från dess ägare!
		-- J. R. R. Tolkien

%
För gin, i grymSober sanning,Levererar bränsletFör flammande ungdom.
		-- Noel Coward

%
För adelskap är inte i bedrifter av krig,När det gäller att kämpa i gräl rätt eller fel,Men i en sak som sanning inte kan skjuta upp:Han borde själv för att kontrollera och stark,Bara för att hålla Mixt med nåd bland:Och inget otalt en riddare borde taMen för en sanning, eller för den gemensamma skull.
		-- Stephen Hawes

%
"Force är men kanske" läraren sa--"Denna definition är bara."Pojken sade intet utan tänkte i stället,Minnas hans dunkade huvudet:"Force är kanske inte men måste!"
		-- Stephen Hawes

%
Fyra vara de saker jag är klokare att veta:Sysslolöshet, sorg, en vän, och en fiende.Fyra vara saker som jag skulle varit bättre utan:Kärlek, nyfikenhet, fräknar, och tvivel.Tre vara de saker jag aldrig uppnå:Avund, innehåll och tillräcklig champagne.Tre vara de saker jag skall ha tills jag dör:Skratt och hopp och en strumpa i ögat.
		-- Dorothy Parker, "Inventory" [or "Not so Deep as a Well"?]

%
Vänner, romare, Hipsters,Låt mig clue du;Jag kommer att lägga ner Caesar, inte att dansa honom.Torget sparkar några katter på vistelse med dem;Höft bitar, som går ner under,så låt den ligga med Caesar. Den svala BrutusGav det meddelande som du: Caesar hade stora ögon;Om det är ljudet, är någon copping en grund,Och, som, gammal Caesar verkligen ställa dem rakt.Här, copacetic med Brutus och tapparna, -för Brutus är en riktigt cool katt;Så är de alla, alla coola katter, -Kommer jag att göra detta spelning på Caesars om.
		-- Dorothy Parker, "Inventory" [or "Not so Deep as a Well"?]

%
Från alltför mycket kärlek att leva,Från hopp och rädsla fri,Vi tackar med kort tacksägelse,Allt vad gudar kan vara,Att inget liv lever för evigt,Att döda män stiga upp aldrig,Att även den weariest floden slingrar någonstans säkert till havs.
		-- Swinburne

%
Komma i kontakt med dina känslor av fientlighet mot den döende ljuset.
		-- Dylan Thomas [paraphrased periphrastically]

%
Ut, din gamla Wight! Försvinna i solljuset!Skrumpnar som kall dimma, som vinden går klagan,Ut i de karga land långt bortom bergen!Kom aldrig hit igen! Lämna din skottkärra tom!Förlorade och glömmas bort, mörkare än mörkret,När portarna står för alltid stänga, tills världen lagade.
		-- J. R. R. Tolkien

%
Gibsons Springtime Song (till tonerna av "Deck the Halls"):'Tis säsongen att jaga mousies (Fa la la la la, la la la la)Rycka dem ur deras små housies (...)Först jaga vi dem "runt fältet (...)Sedan har vi dem för en måltid (...)Slänga dem här och fånga dem där (...)Se dem flyger genom luften (...)Titta på dem flyga och höra dem skrika (...)Fallande möss har stor vädjan (...)Se jägaren sträckt framför oss (...)Han jagade möss i skog och mark (...)Se honom rengöra sina långa vita whiskers (...)Av blodet av lite nötkreatur (...)
		-- J. R. R. Tolkien

%
Gil-Galad var en Elven-kung.Av honom Harpers tyvärr sjunga:den sista vars rike var fria och rättvisamellan bergen och havet.Hans svärd var lång, hans lans var angelägen,hans lysande rodret fjärran sågs;de oräkneliga stjärnorna på himmelen fältåterspeglades i hans silver sköld.Men länge sedan red han bort,och där han bor ingen kan säga;för i mörkret föll hans stjärnai Mordor där skuggor är.
		-- J. R. R. Tolkien

%
Gimme Twinkies, gimme vin,    Gimme jeans av Calvin Kline ...Men om du delar dessa atomer bra,    Mama hålla dem utanför dessa gener av mina!Gimme finnar, ta min deg,    Gimme arsenik i min Jelly Roll ...Ring djävulen och sälja min själ,    Men mamma hålla dem-atomer helhet!
		-- Milo Bloom, "The Split-Atom Blues," in "Bloom County"

%
Ge mig uttalade, upprätt, den manliga fiende,Fet Jag kan möta - kanske kan vända sin slag!Men alla plågor, bra Heaven, din vrede kan skicka,Rädda mig, åh rädda mig från uppriktig vän.
		-- George Canning

%
Ge mig dina elever, dina sekreterare,Dina huddled författare längtan att andas fritt,Eländiga avfall av din Selectric III: s.Ge dessa hemlösa, maskinskriverska-kastade till mig.Jag lyfter min disk bredvid processorn.
		-- Inscription on a Word Processor

%
Gå fridfullt bland buller och avfall,Och kom ihåg vad komfort det kan finnas i att äga en bit därav.Undvik tysta och passiva personer, såvida du inte är i behov av sömn.Rotera dina däck.Tala glowingly av dem är större än dig själv,Och lyssna väl deras råd - trots att de är kalkoner.Vet vad de ska kyssa - och när.Kom ihåg att två fel aldrig göra rätt,Men att tre gör.Där det är möjligt, sätta folk på "HOLD".Tröstas, som med tanke på all torka och besvikelse,Och trots de förändrade öden tid,Det finns alltid en stor framtid i datorn underhåll.Du är en lyckträff av universum ...Du har ingen rätt att vara här.Om du kan höra det eller inte, universumSkrattar bakom ryggen.
		-- National Lampoon, "Deteriorata"

%
Gå fridfullt bland buller och avfall, och kom ihåg vilket värde det kanvara att äga en bit därav.
		-- National Lampoon, "Deteriorata"

%
Gud vila ye CS studenter nu är lagren på trumman borta,Låt inget du bestörtning. Skivan är vinglar också.VAX är nere och kommer inte att vara upp, har vi hittat en bugg i Lisp, och AlgolFram till första maj. Kan inte säga falska ifrån sant.Programmet som berodde detta morgonen, och nu finner vi att vi inte kan fåKommer inte att skjutas upp, säger de. På Berkeleys 4,2.(Kör) (kör)Vi har precis fått ett samtal från december, och nu en del glada nyheter för dig,De skickar utan dröjsmål Nätverkets också död,En bildskärm som kallas RSuX Vi måste skriva ut dina filer påDet tar nio hundra K. radskrivare istället.Personalen begått självmord, handläggningstid är nitton veckor.Vi ska begrava dem i dag. Och bara kort läses.(Kör) (kör)Och nu vill vi säga till dig CHORUS: Åh, budskap om tröst och glädje,Innan vi går bort, komfort och glädje,Vi hoppas de nyheter vi har fört till dig Åh, budskap om tröst och glädje.Kommer inte förstöra hela dagen.Du har ett annat program på grund av, i morgon, förresten.(kör)
		-- to God Rest Ye Merry Gentlemen

%
Gold coast slavskepp på väg till bomullsfältSäljs på en marknad i New OrleansÄrrad gammal slaver vet att han gör alrightHör honom piska kvinnor, precis runt midnattAh, farinsocker hur kommer du smaka så bra?Ah, farinsocker precis som en ung flicka börTrummor som slår kallt engelskt blod går varmLady av huset wonderin "där det kommer att slutaHus pojke vet att han gör alrightDu bör en hörde honom precis runt midnatt....Jag slår vad om din mamma var tält show drottningOch alla hennes väninnor var sweet sixteenJag är ingen skolpojke men jag vet vad jag gillarDu skulle ha hört mig bara runt midnatt.
		-- Rolling Stones, "Brown Sugar"

%
Har fru och barn i Baltimore Jack,Jag gick ut för en åktur och aldrig kom tillbaka.Som en flod som inte vet var det är flytande,Jag tog fel och jag bara fortsatte att gå.Alla har en hungrig hjärta.Alla har en hungrig hjärta.Lägg ner dina pengar och du spelar din del,Alla har en hungrig hjärta.Jag träffade henne i en Kingstown bar,Vi blev kär, jag visste att det skulle sluta.Vi tog vad vi hade och vi slet isär,Nu är jag här nere i Kingstown igen.Alla behöver en plats att vila,Alla vill ha ett hem.Inte göra någon skillnad vad ingen sägerÄr inte ingen gillar att vara ensam.
		-- Bruce Springsteen, "Hungry Heart"

%
Grafik blinda ögon.Ljudfiler deafen örat.Musklick bedöva fingrarna.Heuristik försvagar sinnet.Alternativ vissna hjärtat.The Guru observerar nätetmen litar hans inre syn.Han gör saker att komma och gå.Hans hjärta är så öppet som etern.
		-- Bruce Springsteen, "Hungry Heart"

%
H: Om en "GOBLIN (HOB) waylays dig,Skiva upp honom innan han dödar dig.Ingenting gör att du ser en sluskSom löper från en HOB'LIN (GOB).
		-- The Roguelet's ABC

%
"Hade han och jag men mötteAv några gamla antika inn, men varierade som infanteri,Vi borde ha satt oss ner till våta och stirrar ansikte mot ansikte,Rätt många nipperkin! Jag sköt på honom som han på mig,Och dödade honom i hans ställe.Jag sköt honom död på grund -Eftersom han var min fiende, han trodde att han skulle "lista, kanske,Bara så: min fiende naturligtvis han var; Off-hand som - precis som jag -Det är tillräckligt tydlig; men var utan arbete - hade sålt sina fällorIngen annan anledning varför.Ja; pittoreska och nyfiken krig är!Du skjuter en kollega nerMan skulle kunna behandla, om de uppfylls där någon bar ärEller bidra till en halv krona. "
		-- Thomas Hardy

%
Hälften ett bi, filosofiskt, måste sakens natur halv inte vara.Men halv biet har fått vara, gentemot sin enhet. Se?Men kan ett bi sägas vara eller inte vara en hel bee,När halv biet inte är ett bi, på grund av någon gammal skada?
		-- Thomas Hardy

%
Hängande i tyst desperation är den engelska vägen.
		-- Pink Floyd

%
Papperskopior och ChmodOch alla tror datorer är opersonligakalla diskdrives hårdvaru bildskärmaranvändar fientlig programvaranaturligtvis de är bara bitar och bytesoch tecken och strängaroch filerbara några gamla textfiler från min gamla pojkvänberättade han älskar mig ochhan kommer att ta hand om mighelt enkelt en kasserad utskrift av en väns katalogdjupa intima hemligheter ochhur han inte litar på migkunde inte skada mig mer om de doftande i lavendel eller mögelpå personlig brevpapper
		-- terri@csd4.milw.wisc.edu

%
Hark, Herald Tribune sjunger,Reklam fantastiska saker.Änglar vi har hört på högBerätta att gå ut och köpa.
		-- Tom Lehrer

%
Har du någonsin känt som en sårad kohalvvägs mellan en ugn och en betesmark?går i en trance mot en gravidsjutton-årig hemmafrutvå dagar gamla kokbok?
		-- Richard Brautigan

%
Har du sett hur Sonnys brännande,Liksom några ljusa erotiska stjärna,Han lyser upp målet,Och höjer temperaturen.
		-- The Birthday Party, "Sonny's Burning"

%
Har du sett den gamle mannen i den nedlagda marknaden,Sparka upp tidningarna i sina utslitna skor?I hans ögon du ser ingen stolthet, händer hänga löst på sin sidaGårdagens papper, berättar gårdagens nyheter.Hur kan du säga att du är ensam,Och säga dig solen inte skiner?Låt mig ta dig i handenLeder dig genom gatorna i LondonJag ska visa dig något att få dig att ändra dig ...Har du sett den gamle mannen utanför havs mannens uppdragMinnen blekning liksom de metallbanden som han bär.I vår vinter stad regnet gråter lite syndFör en mer bortglömd hjälte och en värld som inte bryr sig ...
		-- The Birthday Party, "Sonny's Burning"

%
Har du sett den well-to-do, upp och ned Park Avenue?På den berömda huvudgata, med näsan i luften,Höga hattar och Arrow kragar, vita spats och massor av dollar,Spendera varje krona, för en underbar tid ...Om du är blå och du inte vet var du ska gå till,Varför inte gå där mode sitter,...Klädd som en miljon dollar trooper,Försöker hårt för att se ut som Gary Cooper, (super dooper)Kom, låt oss blanda där Rockefeller promenad med stavar,Eller umberellas i sina vantar,Puttin 'on the Ritz....Om du är blå och du inte vet var du ska gå till,Varför inte gå där mode sitter,Puttin 'on the Ritz.Puttin 'on the Ritz.Puttin 'on the Ritz.Puttin 'on the Ritz.
		-- The Birthday Party, "Sonny's Burning"

%
Han hörde att det ofta flygande ljudFötter så lätt som lind-blad,Av musik welling tunnelbana,I dolda håligheter darrande.Nu vissnade lägga odört-skivorna,Och en efter en med suckande ljudViskande föll Beechen bladenI vinter skogsmark vackla.Han sökte henne någonsin, vandra långtNär bladen år var tätt strödda,Med ljus av månen och stråle av stjärnanI frostiga himlen frossa.Hennes mantel glimmade i månen,Som på en kulle-top högt och långtHon dansade, och vid hennes fötter var ströddaEn dimma av silver darrar.När vintern gick, kom hon igen,Och hennes sång släppte plötsligt våren,Liksom stigande lark, och fallande regn,Och smältvatten bubblande.Han såg Elven-blommor vårenOm hennes fötter, och läkt igenHan längtade efter henne att dansa och sjungaVid gräset untroubling.
		-- J. R. R. Tolkien

%
Han trodde att han såg en albatrossDet fladdrade "runt lampan.Han såg igen och såg att det varEn öre frimärke."Du skulle bäst att få hem", sade han,"Nätterna är ganska fuktiga."
		-- J. R. R. Tolkien

%
Den som uppfinner talesätt för andra att ta del avtar längs roddbåt när man går på kryssning.
		-- J. R. R. Tolkien

%
Han som förlorar, vinner loppet,Och parallella linjer möts i rymden.
		-- John Boyd, "Last Starship from Earth"

%
Han har varit som en far för mig,Han är den enda DJ du kan få efter tre,Jag är en all-night musiker i en rock and roll band,Och varför han inte gillar att jag inte förstår.
		-- The Byrds

%
Hennes låser en gammal dam gavHennes kärleksfull mans liv för att rädda;Och män - de hedrade så dame -Vid några stjärnor skänkte hennes namn.Men till vår moderna gift rättvis,Vem skulle ge sina herrar för att rädda sitt hår,Ingen stjärn erkännande har gett.Det finns inte stjärnor tillräckligt i himlen.
		-- The Byrds

%
Här är jag igen precis där jag vet att jag borde inte varaJag har fångats inne i den här fällan för många gångerJag måste ha gått dessa steg och sagt dessa ord entusen gånger innanDet verkar som om jag vet att alla linjer.
		-- David Bromberg, "How Late'll You Play 'Til?"

%
Här sitter jag, förkrossad,Alla inloggade men arbeta Inte startat.Första net.this och net.that,Och en varm smörade bun för net.fat.Chefen kommer förbi, och jag spelar spelet,Då vänder jag tillbaka till net.flame.Finns det ett botemedel (jag behöver era åsikter)För någon instängd i net.news?Jag behöver din hjälp, säger jag mellandäck snyftar,"Orsak kommer jag snart vara införd i net.jobs.
		-- David Bromberg, "How Late'll You Play 'Til?"

%
Här i mitt hjärta, jag är Helen;Jag är Aspasia och Hero, åtminstone.Jag är Judith och Jael och Madame de Sta "el;Jag är Salome, måne i öst.Här i min själ jag Sappho;Lady Hamilton jag, liksom.I mig R 'ecamier tävlar med Kitty O'Shea,Med Dido, och Eva och dålig Nell.Jag är alla de glamorösa damerVid vars vinkande historia skakade.Men du är en man, och ser bara min panna,Så jag stannar hemma med en bok.
		-- Dorothy Parker

%
Här vilar LESTER MOORESHOT 4 gånger med en 0,44NO LESNO MOORE
		-- tombstone, in Tombstone, AZ

%
Hej dol! glad dol! ringa en dong dillo!Ring en dong! hop tillsammans! fal Lal pil!Tom Bom, jolly Tom Tom Bombadillo!
		-- J. R. R. Tolkien

%
Hallå! Kom derry dol! Hop längs mina hearties!Hober! Ponnyer alla! Vi är förtjusta i partier.Låt nu det roliga börjar! Låt oss sjunga tillsammans!
		-- J. R. R. Tolkien

%
Hallå! Kom glatt dol! derry dol! Min älskling!Ljus går väder vind och befjädrade stare.Ner längs enligt Hill, glänsande i solen,Väntar på tröskeln till den kalla starlight,Där min vacker dam är River-kvinnans dotter,Smal som vide-staven, klarare än vattnet.Old Tom Bombadil näckrosor föraKommer hoppande hem igen. Kan du höra honom sjunga?Hallå! Kom glatt dol! derry dol! och glad-oGoldberry, Goldberry, glad gul bär-o!Stackars Willow-man, stoppa du dina rötter bort!Toms bråttom nu. Kväll kommer att följa dag.Tom kommer hem igen näckrosor föra.Hallå! komma derry dol! Kan du höra mig sjunga?
		-- J. R. R. Tolkien

%
Hallå! nu! Kom hoy nu! Vart vill du vandra?Upp, ner, nära eller långt, här, där eller där borta?Sharp-öron, Wise-näsa, Swish-svans och Bumpkin,White-strumpor min lilla pojke, och gamla Fatty Lumpkin!
		-- J. R. R. Tolkien

%
Hej, Hey, Hey spill PDLFör att få lite mer stack;Om detta inte räcker då du förlora alltOch måste pop hela vägen tillbaka.
		-- J. R. R. Tolkien

%
Hickory Dickory Dock,Mössen sprang upp klockan,Klockan slog ett,De andra kom undan med lindriga skador.
		-- J. R. R. Tolkien

%
Hier liegt ein Mann ganz obnegleich;Im Leibe dick, en Suden riket.Wir haben ihn in das Grab gesteckt, Här ligger en man med diverse bristerWeil es uns dunkt ER sei verreckt. Och många synder på huvudet;Vi begravde honom i dag på grund avSåvitt vi kan se, han är död.Sue Bach och skriven av den lokala doggeral catcher;"The Definitive Biografi av PDQ Bach", Peter Schickele
		-- PDQ Bach's epitaph, as requested by his cousin Betty

%
Higgeldy Piggeldy,Hamlet av HelsingörRuggig kritikerna avSläppa bomben:"Phooey på Freud och hanspsyko~~POS=TRUNC -Oidipus Shmoedipus,Jag bara älskar mamma. "
		-- PDQ Bach's epitaph, as requested by his cousin Betty

%
... Hans lärjungar leda honom; han bara gör resten.
		-- The Who, "Tommy"

%
Historien är nyfiken sakerMan skulle kunna tro nu hade vi nogMen faktum kvarstår är jag räddDe gör mer av det varje år.
		-- The Who, "Tommy"

%
Hit dem kex med en annan touch av sås,Bränn att korven bara en match eller två mer gjort.Häll min svarta gamla kaffe längre,Även om det luktar gettin 'starkareEn halv måltid inte nuthin mycket att önska.Låna mig tio, fick jag en feelin 'det ska rädda mig,Med en ornery själ som inte skjuta pool för skojs skull,Om det coat'll passa du wearin,Den Lord'll prise din sharin 'En semi-vän är inte nuthin mycket att önska.Och låt mig halvvägs bli kär,För en del av en ensam natt,Med en halv vacker kvinna i mina armar.Ja, jag kunde halvvägs falla deep--I en snugglin ", lovin hög,Med en halv vacker kvinna i mina armar.
		-- Elroy Blunt

%
Ho! Ho! Ho! till flaskan jag gårAtt läka mitt hjärta och dränka min ve.Regn kan falla och vind kan blåsa,Och många miles fortfarande vara att gå,Men under ett högt träd jag kommer att ligga,Och låt molnen segla förbi.
		-- J. R. R. Tolkien

%
Ho! Tom Bombadil, Tom Bombadillo!Av vatten, trä och berg, genom vass och vide,Genom eld, sol och måne, harken nu och höra oss!Kom, Tom Bombadil, för vårt behov är nära oss!
		-- J. R. R. Tolkien

%
Hop längs mina små vänner, upp Withywindle!Tom händer framåt ljus för att tända.Ner väster sjunker solen; snart kommer du att famlande.När natt skuggor faller, då dörren öppnas,Ut ur winfow-rutor lampan blinkar gult.Fruktar ingen al svart! Lyssna ingen hoary vide!Frukta varken rot eller gren! Tom går innan du.Hej nu! glad dol! Vi kommer att vänta på dig!
		-- J. R. R. Tolkien

%
Hur kan du ha någon pudding om du inte äter ditt kött?
		-- Pink Floyd

%
Hur förtär lilla krokodilFörbättra sitt lysande svans,Och häll vattnet i NilenPå varje gyllene skala!Hur glatt han verkar flina,Hur snyggt sprider klorna,Och välkomnar små fiskar i,Med försiktigt leende käkar!
		-- Lewis Carrol, "Alice in Wonderland"

%
Hur doth VAX s C-kompilatorFörbättra dess objektkod.Och även när vi talar gör detÖka systembelastningen.Hur tålmodigt det verkar köraOch spotta ut felflaggor,Medan användare, med frustration, allaRiv sina kläder till trasor.
		-- Lewis Carrol, "Alice in Wonderland"

%
Dumpty satt på väggen,Humpty Dumpty hade en stor nedgång!Alla kungens hästar,Och alla kungens män,Hade äggröra till frukost igen!
		-- Lewis Carrol, "Alice in Wonderland"

%
Jag kommer alltid att minnas - jag var inte på humör att leka;'Twas ett år sedan November - Jag fick ner min trogna gevärJag gick ut för att skjuta några rådjur och gick ut för att förfölja min byte -På morgonen ljus och tydlig. Vad ett drag jag gjorde den dagen!Jag gick och sköt maximala jag bunden dem till min stötfångare ochSpelet lagar skulle göra det möjligt: ​​Jag körde hem dem på något sätt,Två viltvårdare, sju jägare, två viltvårdare, sju jägare,Och en ko. Och en ko.Lagen var mycket fast, det Folk frågar mig hur jag gör detTog bort mina permit-- Och jag säger, "Det finns inget att det!Den värsta straff jag någonsin fått utstå. Du står bara där lookin söt,Det visar sig att det fanns en anledning. Och när något rör sig, du skjuter "Kor var av säsongen, och Och det finns tio stoppade huvudenEn av jägarna inte var försäkrad. I mitt trofé rum just nu:Två viltvårdare, sju jägare,Och ett renrasigt guernsey ko.
		-- Tom Lehrer, "The Hunting Song"

%
Jag ändra mitt namn till ChryslerJag ska ner till Washington, D.C.Jag kommer att tala om viss makt mäklareVad de gjorde för IacoccaKommer att vara helt acceptabelt för mig!Jag ändra mitt namn till Chrysler,Jag är på väg för den stora mottagande linje.När de lämnar en miljon stor ut,Jag kommer att stå med min hand,Yessir, jag får min!
		-- Tom Lehrer, "The Hunting Song"

%
I B MU B MVi alla B MFör jag B M !!!!
		-- H.A.R.L.I.E.

%
Jag kan leva utanNågon som jag älskarMen inte utanNågon jag behöver.
		-- "Safety"

%
Jag kan se honom a'comin "Med sina stora stövlar på,Med sin stora tummen ur,Han vill få mig.Han vill skada mig.Han vill få ner mig.Men en tid senare,När jag känner mig lite rakare,Jag kommer att stöta en främlingVem kommer att påminna mig om faran,Och då .... jag ska köra honom.Ganska smart för min del!Att hitta min väg ... I mörkret!
		-- Phil Ochs

%
Jag kan inte klaga, men ibland jag fortfarande gör.
		-- Joe Walsh

%
Jag vet inte vad Descartes fick,Men sprit kan göra vad Kant kan inte.
		-- Mike Cross

%
Jag behöver inte några armar runt mig ...Jag behöver inte några droger för att lugna mig ...Jag har sett skriften på väggen.Tro inte att jag behöver något alls.Nej! Tro inte att jag behöver något alls!Allt som allt var det bara tegelstenar i väggen.Allt som allt var det bara tegelstenar i väggen.
		-- Pink Floyd, "Another Brick in the Wall", Part III

%
Jag vill inte argumentera, och jag vill inte slåss,Men det kommer definitivt att vara en part i kväll ...
		-- Pink Floyd, "Another Brick in the Wall", Part III

%
Jag vill inte ha en knipa,Jag vill bara rida på min motorsickle.Och jag vill inte dö,Jag vill bara att rida på min motorcy.Cle.
		-- Arlo Guthrie

%
Jag gav min kärlek en Apple, som inte hade någon kärna;Jag gav min kärlek en byggnad, som inte hade någon golvet;Jag skrev min kärlek ett program, som inte hade någon ände;Jag gav min kärlek en uppgradering, utan cryin ".Hur kan det finnas en Apple, som inte har någon kärna?Hur kan det vara en byggnad, som inte har någon golvet?Hur kan det finnas ett program, som inte har något slut?Hur kan det vara en uppgradering, utan cryin '?En Apples MOS minne använder inte någon kärna!En byggnad som är perfekt, har det ingen brist!Ett program med GOTO, har det inget slut!Jag ljög om uppgraderingen, utan cryin '!
		-- Arlo Guthrie

%
Jag får upp varje morgon, samla mina förstånd.Plocka upp tidningen, läsa obits.Om jag inte är där jag vet att jag är inte död.Så jag äter en bra frukost och gå tillbaka till sängen.Åh, vad vet jag min ungdom är allt använt?Min get-up-and-go har fått upp-och-gick.Men trots allt, jag kan flina,Och tänk på de platser som min utstyrsel har varit.
		-- Pete Seeger

%
Jag hade ett ärende där: samla näckrosor,gröna blad och liljor vita att tillfredsställa min vacker dam,den sista ere årets slut för att hålla dem från vintern,blomma av hennes vackra fötter tills snön smälter.Varje år vid sommarens slut jag gå för att hitta dem för henne,i en bred pool, djup och klar, långt ner Withywindle;där de öppnar först under våren och det de kvar senast.Genom denna pool länge sedan hittade jag floden-dotter,rättvis ung Goldberry sitter i vassen.Söta var hennes sång sedan, och hennes hjärta slog!Och det visade sig vara bra för dig - för nu ska jag inte längregå ner djupt igen längs skogs vatten,nej medan år är gammal. Inte heller ska jag vara passerarOld Man Willow hus denna sida av vår tid,inte förrän den glada våren, när floden-dotterdansar ner withy-väg att bada i vattnet.
		-- J. R. R. Tolkien

%
Jag har en liten skugga som går in och ut med mig,Och vad kan vara användningen av honom är mer än vad jag kan se.Han är mycket, mycket som jag från hälarna upp till huvudet;Och jag ser honom hoppa framför mig, när jag hoppar in i min säng.Det roligaste om honom är hur han gillar att grow--Inte alls som riktiga barn, som alltid är mycket långsam;För han skjuter ibland upp längre, som en Indien-gummiboll,Och han ibland blir så litet att det är ingen av honom alls.
		-- R. L. Stevenson

%
Jag har lärt migAtt stava smårätterSom fortfarande river påVissa människors n'oeuvres.
		-- Warren Knox

%
Jag har massor av saker i mina fickor;Ingen av dem är värt något.Sociopolitiska whines åt sidan,Gan du ger mig, gratis, gratis,Priset på en halv gallonAv Gallo extra dåligOch de flesta av bussresan hem.
		-- Warren Knox

%
Jag tvivlar inte på djävulen flinar,Som hav av bläck jag stänka.Gudar, förlåt min "litterära" sins--Den andra slag spelar ingen roll.
		-- Robert W. Service

%
Jag har den gamla biologiska behov,Jag har den gamla oemotståndliga uppsving,Jag är hungrig.
		-- Robert W. Service

%
Jag visste Leo G. CarrolVar över ett fatNär Tarantula tog till bergen. [ "Slicka det!"]Och jag fick verkligen hetaNär jag såg Jeanette ScottFight en triffid som spottar gift och dödar.Science fiction, dubbel funktionDoktor X kommer att bygga en varelse.Se androider slåss Brad och JanetAnne Francis stjärnor i Forbidden PlanetOh Oh Oh Oh OhVid sent på kvällen, dubbel funktion, bildspel.
		-- The Rocky Horror Picture Show

%
Jag vet inte om du har pratar du gjort sahur förvånad du wuz av levande döda.Du wuz förvånad att de kunde förstå dig ordoch aldrig svara en gång till hela sanningen de hörde.Men inte får fyrkantiga!Det är ingen regel som säger att de fick vård.De kan alltid svär de är döva, stumma och blinda.
		-- The Rocky Horror Picture Show

%
Jag nyligen förlorat en preposition;Det gömde, tänkte jag, under min stolOch ilsket jag ropade, "Perdition!Upp ut ur under där. "Korrektheten är min handbok,Och spretande fraser jag avskyr,Och ändå jag undrade: "Vad skulle han kommaUpp ut ur ramen för? "
		-- Morris Bishop

%
Jag lägger mitt huvud på järnvägsspåren,Waitin för dubbel E.Järnvägen inte köra längre.Dålig dålig ynklig mig. [kör]Dålig dålig ynklig mig, dålig dålig ynklig mig.Dessa unga flickor kommer inte låta mig vara,Herre förbarma dig över mig!Ve mig!Tja, träffade jag en flicka, West Hollywood,Tja, jag inte nämna namn.Men hon verkligen arbetat mig över bra,Hon var precis som Jesse James.Hon arbetade verkligen mig över bra,Hon var en kredit till hennes kön.Hon satte mig igenom några förändringar, pojke,Ungefär som en Waring-blandare. [kör]Jag träffade en tjej på Rainbow Bar,Hon frågade mig om jag skulle slå henne.Hon tog mig tillbaka till Hyatt House,Jag vill inte prata om det. [kör]
		-- Warren Zevon, "Poor Poor Pitiful Me"

%
Jag träffade honom i ett träsk i DagobahOm det bubblar hela tiden som en jätte kolsyrad läskS-O-D-A-sodaJag såg den lilla runt sitter där på en stockJag frågade honom hans namn och i en raspiga röst sade han YodaY-O-D-A Yoda, Yo-Yo-Yo-Yo YodaJo jag har varit runt men jag har aldrig settEn kille som ser ut som en Muppet men han rynkig och gröntOh my Yoda, Yo-Yo-Yo-Yo YodaJag är väl inte dum men jag kan inte förståHur han kan höja mig i luften bara genom att höja sin handOh my Yoda, Yo-Yo-Yo-Yo Yoda, Yo-Yo-Yo-Yo Yoda"Lola" av Kinks
		-- Weird Al Yankovic, "The Star Wars Song," to the tune of

%
Jag måste skapa ett system, eller enslav'd av en annan mans;Jag kommer inte att resonera och jämför; mitt företag är att skapa.
		-- William Blake, "Jerusalem"

%
Jag har aldrig sett en purpurfärgad koJag hoppas att aldrig se enMen jag kan berätta ändåJag skulle hellre se än vara en.Jag har aldrig sett en lila koJag hoppas att aldrig se enMen från mjölken vi får nuDet säkert måste vara enAh, ja, jag skrev "The Purple Cow"Jag är ledsen nu jag skrev detMen jag kan berätta ändåJag ska döda dig om du citerar den.
		-- Gellett Burgess, many years later

%
Jag är skyldig, jag är skyldig,Det är iväg till arbetet jag går ...
		-- Gellett Burgess, many years later

%
Jag hatar verkligen denna förbannade maskinJag önskar att de skulle sälja det.Det gör aldrig riktigt vad jag villMen bara vad jag säger det.
		-- Gellett Burgess, many years later

%
"Jag sa," Preacher, ge mig styrka för runda 5. "Han sade, "Vad du behöver är att växa upp, son."Jag sa, "growin" upp leder till growin gamla,Och sedan dö, och för mig som inte låter som mycket roligt. "
		-- John Cougar, "The Authority Song"

%
Jag såg en man fullfölja Horizon,"Runt, runt de accelererade.Jag stördes på detta,Jag tilltalade mannen,"Det är meningslöst", sa jag."Du kan never--""Du ljuger!" Han grät,och sprang vidare.
		-- Stephen Crane

%
Jag ser en dålig moon rising.Jag ser problem på vägen.Jag ser jordbävningar och Lightnin 'Jag ser dåliga tider idag.Inte att gå runt i kväll,Det är skyldig att ta ditt liv.Det är en dålig månen på uppgång.
		-- J. C. Fogerty, "Bad Moon Rising"

%
Jag ser egenvärdet i ditt öga,Jag hör anbuds tensor i din suck.Bernoulli skulle ha nöjt sig med att döHade han men kända sådana _ a-squared cos 2 (phi)!
		-- Stanislaw Lem, "Cyberiad"

%
Jag skickade ett brev till fisken, sa jag det mycket högt och tydligt,Jag sa till dem, "Detta är vad jag vill." Jag gick och ropade i hans öra.De små fiskarna i havet, men han var mycket hård och stolt,De skickade ett svar tillbaka till mig. Han sa "Du behöver inte skrika så högt."De små fiskarna "svar var och han var mycket stolt och hård,"Vi kan inte göra det, sir, eftersom ..." Han sa "Jag ska gå och väcka dem om ..."Jag skickade ett brev tillbaka att säga att jag tog en vattenkokare från hyllan,Det vore bättre att lyda. Jag gick för att väcka upp dem själv.Men någon kom till mig och sa men när jag fann dörren var låst"De små fiskarna är i sängen." Jag drog och knuffade och sparkade ochknackade,Jag sade till honom, och jag sa att det klart och när jag fann dörren stängdes,"Då måste du väcka dem upp igen." Jag försökte vrida handtaget, men ...	"Är det allt?" frågade Alice.	"Det är allt." sade Humpty Dumpty. "Adjö."
		-- Stanislaw Lem, "Cyberiad"

%
Jag skickade ett meddelande till en annan tid,Men allteftersom dagarna varva ned - detta jag bara kan inte tro,Jag skickade ett meddelande till en annan planet,Kanske är det ett spel - men det jag bara inte kan föreställa sig....Jag träffade någon som tittar på väldigt lik dig,Hon gör det du gör, men hon är en IBM.Hon är endast programmerad att vara mycket trevligt,Men hon är så kall som is, när jag får för nära,Hon berättar att hon gillar mig väldigt mycket,Men när jag försöker röra, hon gör det alltför tydligt....Jag inser att det måste verka så konstigt,Den tiden har omfördelat, men tiden har sista ordet,Hon vet att jag tänker på dig, hon läser mitt sinne,Hon försöker vara ovänlig, hon vet ingenting om vår värld.
		-- ELO, "Yours Truly, 2095"

%
Jag sköt en fråga till nätet.Jag har inte fått något svar ännu, kallas A postat meddelande mig ruttnaMen sju personer gav mig fan för att ignorera mail jag hade aldrig fått;Och sa att jag borde lära sig att stava; En arg budskap frågade mig, VänligenSkicka inte ett sådant dravel utomlands;En advokat skickade mig privat postOch svor att han skulle smälla min röv i fängelse - En netter trodde att det var en bluff:Jag hade nämnt Un * x i min pärla "Livet, lägga till nettopunkt skämt!";Och misslyckades med att lägga till T och M; En annan ringde min grammatik vileOch kritiserade min handstil.Varje dag scanna I varje ämnesradI hopp ämnet blir min;Jag sköt en fråga till nätet.Jag har inte fått något svar ännu ...
		-- Ed Nather

%
Jag stod i framkant,Den östra kusten vid mina fötter."Hoppa!" sade Yoko OnoJag är för rädd och snygg, ropade jag.Gå vidare och ge det ett försök,Varför förlänga plågan måste alla män dö.
		-- Roger Waters, "The Pros and Cons of Hitchhiking"

%
Jag tror att jag aldrig skall höraEn dikt vackrare än öl.De saker som Joes Bar har i omgångar,Med gyllene bas och snöiga locket.De saker som jag kan dricka hela dagenTills min mem'ry smälter bort.Dikter görs av dårar, jag är räddMen bara Schlitz kan göra en öl.
		-- Roger Waters, "The Pros and Cons of Hitchhiking"

%
Jag tror att jag aldrig får seEn skylt vacker som ett träd.I själva verket, om inte skyltar fallerJag kommer aldrig att se ett träd alls.
		-- Ogden Nash

%
Jag tror att jag aldrig får seEn sak så vacker som ett träd.Men som du ser träden har gåttDe gick i morse med gryningen.En loggning firma ut ur stadenKom och hackade träden allt ned.Men jag kommer att lura de smutsiga skunkarOch skriva en helt ny dikt som heter "Trunks".
		-- Ogden Nash

%
"Jag trodde att du sa att du var 20 år gammal!""Som en programmerare, ja", svarade hon,"Och du påstod sig vara mycket nära två meter hög!""Du sa att du var blond, men du ljög!"Åh, hon var en hacker och han var en också,De hade så mycket gemensamt, skulle man kunna säga.De utbytte skämt och dikter, och smarta nya hacka,Och uppmaningar som var söt eller risque ".Han skickade henne en bild av hans bror Sam,Hon skickade ett från vissa tidigare high school dag,Och det kunde ha gått på för resten av livet,Om de inte hade träffat i L.A."Din skägg är en armhåla", sade hon i avsmak.Han svarade: "Din armhålan är ett skägg!"Och de chorused: "Jag tror att jag kunde stå alla de övrigaOm du inte var så helt konstigt! "Om hon inte hade sagt vad han ville höra,Och han hade inte gjort precis samma sak,De skulle ha varit mycket mer ärlig, och aldrig har träffat,Och skulle inte ha haft kul med spelet.		E-post"
		-- Judith Schrier, "Face to Face After Six Months of

%
Jag brukade vara en sådan söt söt sak, 'til de fick tag i mig,Jag öppnade dörrar för gamla damer, jag hjälpte den blinde att se,Jag fick inga vänner "sak de läser tidningarna, de kan inte ses,Med mig, och jag är feelin 'riktiga skott ner,Och jag, eh, feelin "betyder,Inget mer, Mr. Nice Guy,Inget mer, Mr Clean,Inget mer, Mr. Nice Guy,De säger "Han är sjuk, han är oanständigt".Min hund bet mig på benet i dag, min katt klöste mina ögon,Ma kastats ut ur den sociala krets, och pappa har att dölja,Jag gick till kyrkan, inkognito, när alla steg,Pastor Smithy, erkände han mig,Och slog mig i näsan, sade han,(kör)Han sa "Du är sjuk, du är oanständigt".
		-- Alice Cooper, "No More Mr. Nice Guy"

%
Jag föddes i ett fat slaktare knivarTrouble jag älskar och fred jag föraktarVilda hästar sparkade mig i min sidaDå en skallerorm bet mig och han gick bort och dog.
		-- Bo Diddley

%
Jag var eatin "några chop suey,Med en dam i St. Louie,När det plötsligt kommer en knockin på dörren.Och det kläpp, säger han, "Älskling,Rulla rocker ut några pengar,Eller din pappa skjuter en BOV på golvet. "
		-- Mr. Miggle

%
Jag gick hem med en servitris,Som jag alltid gör.Hur jag skulle jag veta?Hon var med ryssarna också.Jag var spelande i Havanna,Jag tog en liten risk.Skicka advokater, vapen, och pengar,Pappa, får mig ut ur denna.
		-- Warren Zevon, "Lawyers, Guns and Money"

%
Jag gick över till min vän, han eatin "en knipa.Jag sa "Hej, vad är happenin '?"Han sade "Nothin '."Försök att sjunga den här låten med den typen av entusiasm;Som om du bara kläm en polis.
		-- Arlo Guthrie, "Motorcycle Song"

%
Jag kommer inte att spela på dragkamp.Jag skulle hellre spela på kram o krig,Där alla kramarIstället för bogserbåtar,Där alla fnittrarOch rullar på matta,Där alla kysser,Och alla grinar,Och alla OmfamningarOch alla vinner.
		-- Shel Silverstein, "Hug o' War"

%
Jag vaknade upp en feelin 'betydergick ner för att spela spelautomatenhjulen vände,och bokstäverna läsa"Bättre gå tillbaka till Tennessee Jed"
		-- Grateful Dead

%
jag skulle vilja vetaVad jag stängsel iOch vad jag stängsel ut.
		-- Robert Frost

%
Jag skulle aldrig gråta om jag hittadeEn blåval i min soppa ...Inte heller skulle jag emot ett piggsvinInuti ett hönshus.Ja livet är bra när saker kombinera,Som skinka nötkött chow mein ...Men herre, den här gången tror jag att jag har något emot,De har lagt syra i min regn.
		-- - Milo Bloom

%
Jag skulle hellre skrattar med syndare,Än gråta med de heliga,Syndare är mycket roligare!
		-- Billy Joel, "Only The Good Die Young"

%
Jag ska ge dig direktåtkomst till mitt hjärta,Thoul't berätta alla konstanterna din kärlek;Och så vi två skall alla kärlekens lemman bevisaOch i vår bundna partition aldrig del.Avbryt mig inte - för vad då skall förbli?Abskissan vissa mantissorna, moduler, lägen,En rot eller två, en torus och en nod:Inversen av min vers, en noll domän.Jag ser egenvärdet i ditt öga,Jag hör anbuds tensor i din suck.Bernoulli skulle ha nöjt sig med att döHade han men kända sådana a-kvadrat cos 2 (thi)!
		-- Stanislaw Lem, "Cyberiad"

%
Jag ska lära sig spela saxofon,Jag spelar bara vad jag känner.Dricka skotsk whisky hela natten lång,Och dör bakom ratten.De fick ett namn för vinnarna i världen,Jag vill ha ett namn när jag förlorar.De kallar Alabama Crimson Tide,Kalla mig Deacon Blues.
		-- Becker and Fagan, "Deacon Blues"

%
Jag ser dig ... på den mörka sidan av månen ...
		-- Pink Floyd

%
Jag är en konstnär.Men det är inte vad jag verkligen vill göra.Vad jag verkligen vill göra är att vara en sko försäljare.Jag vet vad du ska säga -"Dreamer Få huvudet ur molnen."Okej! Men det är vad jag vill göra.Istället måste jag gå på att måla hela dagen lång.Världen borde göra en plats för sko försäljare.
		-- J. Feiffer

%
Jag är fri - och frihet smakar av verkligheten.
		-- The Who

%
Jag är lika tråkigt som tråkigt kan vara!Jag har saknat din speciella datum.Säg att du inte är arg på migMin deklaration är sent.
		-- Modern Lines for Modern Greeting Cards

%
jag lever så långt bortom min inkomst som vi nästan kan sägas varalever åtskilda.
		-- e. e. cummings

%
Jag är N-ari trädet, jag,N-ari trädet, jag, jag.Jag får genomkorsas av tolken intill,Hon genomkorsas mig sju gånger tidigare.Och ev'ry gången var det en N-faldig (N-ary!)Aldrig skulle aldrig göra en binär. (Nej herrn!)Jag är 'er åttonde träd som var N-ary.N-ari trädet jag, jag,N-ari trädet jag.
		-- Stolen from Herman's Hermits

%
Jag är så olycklig utan dig det är nästan som att ha dig härHon fick guldgruva, fick jag ShaftNär My Love kommer tillbaka från damrummet Kommer jag vara för gammal för att bry sig?Jag vet inte om att ta livet av mig eller bowlaDrop Kick Me, Jesus, genom målstolparna of Life
		-- Unattributed song title.

%
Jag är väldigt bra på integral och differentialkalkyl,Jag vet de vetenskapliga namnen på varelser animalculous;Kort sagt, i frågor växt-, djur- och mineral,Jag är mycket modell av en modern generalmajor.
		-- Gilbert & Sullivan, "Pirates of Penzance"

%
Jag har varit på denna ensamma väg så länge,Är det någon som vet om det går,Jag minns förra gången tecknen pekade hem,En månad sedan.
		-- Carpenters, "Road Ode"

%
Jag har byggt en bättre modell än den i Data GeneralFör databaser växt-, djur- och mineralMin OS hanterar processorer med multiplexerade dualitet;Min PL / 1 kompilatorn visar imponerande funktionalitet.Min lagringssystem är bättre än magnetisk kärna polaritet,Du behöver aldrig bry checkar ut en bit för paritet;Det finns inte någon anledning att installera icke-statiska golv mattor;Min hårddisk har kapacitet för rörlig formatering.Jag känner mig tvungen att tala om vad jag vet är en skadeglad punkt:Det finns gott om plats i minnet för variabler floating-point,Vilket visar för inmatning växt-, djur- och mineralJag har byggt en bättre modell än den i Data General."Modern Generalmajor", från "Pirates of Penzance"av Gilbert & Sullivan)
		-- Steve Levine, "A Computer Song" (To the tune of

%
Jag har äntligen hittat den perfekta tjejen,Jag kunde inte begära mer,Hon är döv och stum och överkönsbestämmas,Och äger en spritbutik.
		-- Steve Levine, "A Computer Song" (To the tune of

%
I / O, I / O,Bär det av till disk I går,Lite eller byte för att läsa eller skriva,I / O, I / O, I / O ...
		-- Steve Levine, "A Computer Song" (To the tune of

%
jagärintemycketlyckligverkandenöjdnärhelstframträdandevetenskapsmänovermagnifyintellektuellupplysning
		-- Steve Levine, "A Computer Song" (To the tune of

%
IBM hade en PL / I,Dess syntax värre än JOSS;Och överallt detta språk gick,Det var en total förlust.
		-- Steve Levine, "A Computer Song" (To the tune of

%
Om en nation förväntar att vara okunnig och fri,... Förväntar sig det som aldrig var och aldrig kommer att bli.
		-- Thomas Jefferson

%
Om ett system administreras klokt,användarna kommer att nöja.De tycker hacka sin kodoch inte slösa tid att genomföraarbetsbesparande skalskript.Eftersom de innerligt älskar sina kontonDe är inte intresserade av andra maskiner.Det kan finnas telnet, rlogin, och ftp,men dessa inte åt några värdar.Det kan finnas en arsenal av sprickor och skadlig kod,men ingen någonsin använder dem.Folk tycker om att läsa sin e-post,ta nöje i att vara med sina diskussionsgrupper,spendera helger arbetar på deras terminaler,glädje i förehavanden på platsen.Och även om nästa systemet är så näraatt användarna kan höra sina viktigaste klick och Biff piper,de är nöjda med att dö av ålderdomutan att någonsin ha gått att se det.
		-- Thomas Jefferson

%
Om allt är sant att jag tror,Det finnas fem skäl till varför man bör dricka;Goda vänner, gott vin, eller vara torr,Eller så att vi bör vara med-och-av,Eller någon annan anledning varför.
		-- Thomas Jefferson

%
Om alla hav var bläck,Och alla vassen var pennor,Och alla himlen var pergament,Och alla män kunde skriva,Dessa skulle inte räckaAtt skriva ner alla byråkratiAv denna regering.
		-- Thomas Jefferson

%
Om en S och en I och ett O och ett UMed ett X i slutet stava Su;Och ett E och en Y och en E stavnings I,Be vad är en speller att göra?Då, om också en S och en I och en GOch en hed stavningssidan,Det finns inte mycket kvar för en stavningskontroll att göraMen att gå begå siouxeyesighed.
		-- Charles Follen Adams, "An Orthographic Lament"

%
Om Dr Seuss Var en teknisk skribent .....Här är ett enkelt spel att spela.Här är en lätt sak att säga:Om ett paket träffar en ficka på ett uttag på en port,Och bussen avbryts som en sista utväg,Och adressen till minnet gör din diskett avbryta,Då uttaget paket fickan har ett fel att rapportera!Om markören hittar ett menyalternativ, följt av ett streck,Och ikonen dubbelklicka sätter ditt fönster i papperskorgen,Och dina data är skadad "orsak indexet inte hash,då din situation är hopplös, och systemets gonna krascha!Du kan inte säga det? Vad synd, sir!Vi hittar du ett annat spel, sir.Om etiketten på kabeln på bordet på ditt hus,Säger nätverket är anslutet till knappen på musen,Men dina paket vill tunneln på ett annat protokoll,Det är flera gånger avvisats av skrivaren ner i korridoren,Och skärmen är alla snedvrids av biverkningar av Gauss,Så dina ikoner i fönstret är vågiga som en blöta,Då kan man lika gärna starta och gå ut med en smäll,"Orsaka så säker som jag är en poet, sucker gonna hänga!När en kopia av din diskett blir slarvigt på disken,Och mikrokoden instruktionerna orsaka onödig RISCDå måste man blinka ditt minne och du vill att ramma din rom.Snabbt stänga av datorn och se till att berätta för din mamma!
		-- DementDJ@ccip.perkin-elmer.com (DementDJ) [rec.humor.funny]

%
Om jag kunde läsa ditt sinne, kärlek,Vilken berättelse dina tankar kunde berätta,Precis som en häftad roman,Den typ apoteket säljer,När du når den delen där de sorger kommer,Hjälten skulle vara mig,Hjältar misslyckas ofta,Du kommer inte att läsa den där boken igen, eftersomslutet är alldeles för svårt att ta.Jag går bort, som en filmstjärna,Vem får brännas i en trevägs-skript,Ange nummer två,En film drottningen att spela scenenAtt föra ut allt det goda i mig,Men nu, kärlek, låt oss vara verkligtJag trodde aldrig att jag skulle kunna agera på detta sätt,Och jag måste säga att jag bara inte få det,Jag vet inte var vi gick fel men känslan är bortaOch jag bara inte kan få tillbaka ...
		-- Gordon Lightfoot, "If You Could Read My Mind"

%
Om jag kunde hålla min penna i mitt hjärta,Jag skulle spilla det hela scenen.Skulle det tillfredsställa dig, skulle den glida på genom ya,Skulle du tror att pojken var konstigt?Är han inte konstigt?...Om jag kunde sticka en kniv i mitt hjärta,Självmord höger på scenen,Skulle det vara tillräckligt för din tonåring lust,Skulle det hjälpa att lindra smärtan?Ease din hjärna?
		-- Rolling Stones, "It's Only Rock'N Roll"

%
Om jag inte köra runt parken,Jag är ganska säker på att göra min markering.Om jag i sängen varje natt med tio,Jag kan få tillbaka mitt utseende igen.Om jag avstå från kul och sådant,Jag kommer förmodligen att uppgå till mycket;Men jag ska stanna som jag är,Eftersom jag inte ett dugg.
		-- Dorothy Parker

%
Om jag lovade dig månen och stjärnorna, skulle du tro det?
		-- Alan Parsons Project

%
Om jag reste till slutet av regnbågenSom Dame Fortune hade för avsikt,Murphy skulle vara där för att berättaPotten är i andra änden.
		-- Bert Whitney

%
Om forskarna författade barnvisor ...Little Miss Muffet satt på hennes glutealregionen,Äta komponenter av syrad mjölk.Vid minst ett tillfälle,längs kom en spindeldjur och satte sig bredvid henne,Eller åtminstone i sin närhet,Och fick henne att känna en överväldigande, men inte förlamande, rädsla,Som motiverade patienten att lämna området ganska snabbt.
		-- Ann Melugin Williams

%
Om hon inte hade varit koppar i sina joner,Hennes form ovoidal,Deras romans kan ha blomstrade.Men han byggde tetraedrisk i sin form,Hans joner järn,Kärlek kan inte låta bli att dö,Uncatylised, inert, och undernärd.
		-- Ann Melugin Williams

%
Om du hade bara en minut att andas,Och de gav er en sista önskan,Vill du be om någotSom en annan chans?
		-- Traffic, "The Low Spark of High Heeled Boys"

%
Om du håller ett lager av sprit i ditt skåp,Det är smart att hålla ett lås på ditt lager.Eller någon joker som är slicker,Kommer lura dig om din sprit,Om du misslyckas med att låsa din sprit med ett lås.
		-- Traffic, "The Low Spark of High Heeled Boys"

%
Om du är orolig av jordbävningar och kärnvapenkrig,Samt av trafik och brott,Överväga hur bekymmersfri gophers ärÄven lever på grävt tid.
		-- Richard Armour, WSJ, 11/7/83

%
Il brilgue: les t ^ Oves libricilleuxSe gyrent et frillant dans le guave,ENM ^ im 'es sont les gougebosquex,Et le m ^ omerade horgrave.Es Brilig krig. Die Schlichte TovenWirrten und wimmelten i Waben;Und aller-mumsige BurggovenDir mohmen Rath ausgraben.
		-- Lewis Carrol, "Through the Looking Glass"

%
In / användare3 gjorde Kubla KahnEn ståtlig nöje kupol dekret,Var / bin, sprang den heliga flodenGenom Test Suites measureless till ManNer till en Brun C.
		-- Lewis Carrol, "Through the Looking Glass"

%
I varje jobb som måste göras, det finns ett inslag av nöje.Hitta det roliga och knäpp! Jobbet är ett spel.Och varje uppgift du göra, blir en bit av kakan,en lärka, en spree; Det är mycket tydligt att se.
		-- Mary Poppins

%
I gymnasiet i BrooklynJag var baseball manager,stolt som jag kunde varaJag jagade baseballs,samlats kastas fladdermössdelade ut handdukar småningom köpte jag min egenDet var mycket viktigt arbete, men det var mörkblå medanför en liten spastisk unge, de officiella var grönmen jag var en teammedlem Ingen har någonsin sagt någotNär laget fick med mig om min blå jacka;deras uppvärmning jackor killarna var mina vännerJag fick inte en Ändå skada mig hela åretEndast den vanliga laget att bära den blå jackafick dessa jackor, och bland alla dessa grönasäkert inte en chef Redan nu fyrtio år efter,Jag minns fortfarande den där jackanoch minnet går på skada.
		-- Bart Lanier Safford III, "An Obscured Radiance"

%
I Riemann, Hilbert eller i BanachrumLåt upphöjd och nedsänkt går deras väg.Våra asymptoter inte längre ur fas,Vi ska möta, räkna, ansikte mot ansikte.
		-- Stanislaw Lem, "Cyberiad"

%
I dimestores och busstationerFolk talar om situationerLästa böcker upprepa citatDra slutsatser på väggen.
		-- Bob Dylan

%
Tidigt på morgonen kön,Med en notering i min hand.Med ett bekymmer i mitt hjärta, det på terminal nummer 9,Waitin 'här i Ceras-land. Pascal kör redo att gå.Jag är en lång väg från vila, men jag Waitin i kön,Hur jag saknar en god måltid så. Med denna kod som någonsin växer.I början av mornin kö, nu lobbyn stolar är mjuka,Med ingen plats att gå. Men det kan inte göra kön agera snabbt.Hej, där det går min vän,Jag har flyttat upp en äntligen.Morning Rain "av G. Lightfoot
		-- Ernest Adams, "Early Morning Queue", to "Early

%
I landet av mörkret Ship avSun drivs av Grateful Dead.
		-- Egyptian Book of the Dead

%
I denna dalSlit och syndHuvudet växer skalligMen inte hakan.
		-- Burma Shave

%
I Xanadu gjorde Kubla KhanEn ståtlig nöje kupol kungörelse:Där Alph, den heliga floden, sprangGenom bergrum omätliga för människanNer till en sunless hav.Så två gånger fem miles från grogrundMed murar och torn var gördlad runt:Och det fanns trädgårdar ljus med slingrande rännilar,Där blommade många en rökelse bärande träd;Och här var skog gamla som gatan,Omsluter soliga platser av grönska.
		-- S. T. Coleridge, "Kubla Kahn"

%
I Xanadu gjorde Kubla Khan ett stately nöje kupol kungörelseMen bara om NFL till en franchise skulle hålla.
		-- S. T. Coleridge, "Kubla Kahn"

%
Till kärlek och ut igen,Således gick jag och därför går jag.Skona din röst, och hålla pennan:Väl och bittert vet jagAlla låtar någonsin sjungit,Alla ord någonsin sagt;Kan det vara så, när jag var ung,Någon tappade mig på mitt huvud?
		-- Dorothy Parker, "Theory"

%
Det kan inte ses, inte kan kännas,Kan inte höras, inte kan smälta.Det ligger bakom startar och under kullar,Och tomma hål fyller.Det kommer först och följer efter,Slutar liv, dödar skratt.
		-- Dorothy Parker, "Theory"

%
Det hänger ner från ljuskronaIngen vet riktigt vad det görDess färg är udda och dess form är konstigtDet avger en högtravande surrDen växer ett par fötter varje dagoch slingrar med slags en ryckningInget fel det orsaka det kommer frånen besökande farbror som är rik!
		-- To "It Came Upon A Midnight Clear"

%
Det hände för länge sedanI den nya magiskt landIndianerna och buffelExisterade hand i handIndianerna behövde matDe behöver skinn till ett takDe tog bara vad de behövdeOch buffel sprang lösMen sedan kom den vite mannenMed sin tjocka och tomt huvudHan kunde inte se förbi sin plånbokHan ville alla buffalo dödaDet var tråkigt, ack så tråkigt.
		-- Ted Nugent, "The Great White Buffalo"

%
Det är inte bra för en människa att vara utan kunskap,och den som gör brådska med fötterna saknar sin väg.
		-- Proverbs 19:2

%
Det brukade vara roligt var iAvskiljning och döda.På ett annat ställe och tidJag gjorde det för spänning.
		-- Lust to Love

%
Det var en gång för mycketEtt ord för fåDet var allt för mycket för mig och digDet fanns en väg att gåInget mer vi kunde göraEn gång för mångaEtt ord för få
		-- Meredith Tanner

%
Det är snabbare hästar,Yngre kvinnor,Äldre whisky ochMer pengar.
		-- Tom T. Hall, "The Secret of Life"

%
Det kommer att bli bra,Det är nästan midnatt,Och jag har två flaskor vin.
		-- Tom T. Hall, "The Secret of Life"

%
Det är bara ett hopp till vänsterOch sedan ett steg åt höger.Sätt händerna på höfternaOch dra knäna i tät.Det är bäcken dragkraftDet blir verkligen du insa-a-a-a-aneLåt oss göra tidsförskjutning IGEN!
		-- Rocky Horror Picture Show

%
Det är bara hyreshus regler,Så allt du 'utrymmet hus dårarKom ihåg: en mans taket är en annan mans golv.En mans taket är en annan mans golv.
		-- Paul Simon, "One Man's Ceiling Is Another Man's Floor"

%
Det är så härÄven samurajhar nallar,och även nallarbli full.
		-- Paul Simon, "One Man's Ceiling Is Another Man's Floor"

%
Det är inte mot någon religion att vilja göra sig av med en duva.
		-- Tom Lehrer, "Poisoning Pigeons in the Park"

%
Det är så förvirrande att välja sida i stundens hetta,bara för att se om det är riktigt,Oooh, det är så erotisk har du berätta hur det ska kännas,Men jag undvika alla hårda kalla fakta som jag fick att möta,Så fråga mig bara en fråga när denna magiska natten är igenom,Kan det ha varit vem som helst eller gjorde det måste vara du?
		-- Billy Joel, "Glass Houses"

%
John Dame maj OscarVar homosexuell var Whitty Var WildeMen Gerard Hopkins men John Greenleaf men ThorntonAdes Manley Var Whittier Var Wilder
		-- Willard Espy

%
Johannes Döparen efter förgiftning en tjuv,Tittar upp på sin hjälte, Commander-in-Chief,Säger berätta stor ledare, men se det kortFinns det ett hål för mig att bli sjuk i?Commander-in-Chief svarar honom samtidigt som jagar en fluga,Säger död till alla dem som skulle gnälla och gråta.Och släppa en skivstång han pekar mot himlen,Att säga solen är inte gult, det är kyckling.
		-- Bob Dylan, "Tombstone Blues"

%
Bara en låt innan jag går, går igenom säkerhetskontrollenTill den det berör, höll jag henne så länge.Reser två gånger ljudets hastighet Hon såg slutligen på mig kär,Det är lätt att bli bränd. Och hon var borta.När visar var över bara en låt innan jag går,Vi var tvungna att komma tillbaka hem till en lektion läras.Och när vi öppnade upp dörren Reser två gånger ljudets hastighetJag var tvungen att vara ensam. Det är lätt att bli bränd.Hon hjälpte mig med min resväska,Hon står framför mina ögon,Driver mig till flygplatsenOch till den vänliga skies.
		-- Crosby, Stills, Nash, "Just a Song Before I Go"

%
Bara maskiner att göra stora beslut,Programmeras av män för medkänsla och vision,Vi kommer att vara ren när deras arbete är gjort,Vi kommer att vara evigt fri, ja, evigt ung,Vad en vacker värld kommer detta att vara,Vilken härlig tid att vara fri.
		-- Donald Fagon, "What A Beautiful World"

%
`Bara plats för en Snark!" Bellman ropade,När han landade hans besättning med omsorg;Stöd varje människa på toppen av tidvattnetAv ett finger sammanflätade i håret."Bara plats för en Snark! Jag har sagt det två gånger:Som ensam bör uppmuntra besättningen.Bara plats för en Snark! Jag har sagt det tre gånger:Vad jag berätta tre gånger är sant. "
		-- Donald Fagon, "What A Beautiful World"

%
`Bara plats för en Snark!" Bellman ropade,När han landade hans besättning med omsorg;Stöd varje människa på toppen av tidvattnetAv ett finger sammanflätade i håret.`Bara plats för en Snark! Jag har sagt det två gånger:Som ensam bör uppmuntra besättningen.Bara plats för en Snark! Jag har sagt det tre gånger:Vad jag berätta tre gånger är sant. "
		-- Donald Fagon, "What A Beautiful World"

%
Bara går morse, låt de mig att du var borta,Suzanne, planer de gjort sätta stopp för dig,Jag gick ut i morse och jag skrev ner den här låten,Bara inte kan komma ihåg vem du ska skicka det till ...Åh, jag har sett eld och jag har sett regn,Jag har sett soliga dagar som jag trodde skulle aldrig slut,Jag har sett ensamma gånger när jag inte kunde hitta en vän,Men jag har alltid trott att jag skulle se dig igen.Trodde jag skulle se dig en gång igen.
		-- James Taylor, "Fire and Rain"

%
K: Cobalt metall, hård och glänsande;Cobol s ordrik och innestängande;Kobolds störta när du slår dem;Inte mår dåligt, är det svårt att tycka om dem.
		-- The Roguelet's ABC

%
Håll gamla länder, din storied pompa! gråter honMed tysta läppar. Ge mig era trötta, era fattiga,Din hopkrupen massorna längtan att andas fritt,Eländiga avfall av din myllrande stranden.Överför dessa, hemlösa, storm-kastade mig ...
		-- Emma Lazarus, "The New Colossus"

%
Knock Knock ... (vem är det?) Eter! (Eter vem?) Eter kanin ... Ja![kör]Yeay!Bo på Happy sidan, alltid på den lyckliga sidan,Bo på Happy sidan av livet!Bum bum bum bum bum bumDu kommer att känna någon smärta, som vi kör du galen,Så Bo på Happy sidan av livet!Knock Knock ... (vem är det?) Anna! (Anna vem?)En annan eter kanin ... [chorus]Knock Knock ... (vem är det?) Stilla! (Stilla vem?)Ytterligare en annan eter kanin ... [chorus]Knock Knock ... (vem är det?) Yetta! (Yetta vem?)Ännu en eter kanin ... [chorus]Knock Knock ... (vem är det?) Cargo! (Last vem?)Cargo beep beep och köra över eter kanin ... [chorus]Knock Knock ... (vem är det?) Bu! (Boo vem?)Gråt inte! Eter kanin vara tillbaka nästa år! [kör]
		-- Emma Lazarus, "The New Colossus"

%
Mina damer och herrar, Hobos och Tramps,Skelögd myggor och bowlegged myror,Jag kommer innan du att stå bakom digBerätta om något som jag inte vet någonting om.Nästa torsdag (vilket är bra fredag),Det kommer att finnas en konvention som hölls iKvinnors Club som är strikt för Män.Inträdet är gratis, betala på dörren,Dra upp en stol och sitta på golvet.Det var en sommardag på vintern,Och snön regnar snabbt,Som en barfota pojke med skor på,Stod sitter i gräset.Åh, det ljusa dagen i mitt i natten,Två döda män fick upp till kamp.Tre blinda män att se rent spel,Fyrtio mutes att skrika "Hurra!"Rygg mot rygg, inför de varandra,Drogo sina svärd och sköt varandra.En döv polis hörde buller,Kom och grep de två döda pojkar.
		-- Emma Lazarus, "The New Colossus"

%
Skänkar och Jellyspoons!Jag kommer innan du att stå bakom dig,Berätta något jag inte vet någonting om.Eftersom nästa torsdag kommer att bli långfredagen,Det kommer att finnas en fäder möte, endast mödrar.Bär dina bästa kläder, om du inte har någon,Och snälla stanna hemma om du eventuellt kan vara där.Inträdet är gratis, vänligen betala vid dörren.Har en plats på mig: Vänligen sitta på golvet.Oavsett var du lyckas sitta,Mannen på balkongen kommer säkert spotta.Vi tackar för din ovänlig uppmärksamhet,Och vill nu presentera vår nästa handling:"de fyra hörnen av det runda bordet."
		-- Emma Lazarus, "The New Colossus"

%
Lady, dam, bör du möterEn vars vägar är alla diskret,En som mumlar att hans fruÄr ledstjärna för sitt liv,En som håller försäkra erAtt han var aldrig sant,Aldrig älskat en annan ...Lady, dam, bättre köra!
		-- Dorothy Parker, "Social Note"

%
Nyckelpiga, nyckelpiga,Titta på din akter!Ditt hus brinner,Dina barn kommer att bränna!Så hoppa ni och sjunga, förDen allra första gångenDe fyra linjerna ovanförHar tagits i rim.
		-- Walt Kelly

%
I går kväll träffade jag på trappanEn liten man som inte var där.Han var inte där idag igen.Gee hur jag önskar att han skulle gå bort!
		-- Walt Kelly

%
Latin är ett språk,Död som kan vara.Först dödade romarna,Och nu är det dödar mig.
		-- Walt Kelly

%
Låt mig inte äktenskapet sanna sinnenMedge hinder. Kärlek är inte kärlekSom förändrar när det förändring finnerEller böjar med remover för att ta bort:O, nej! det är en ständigt fast märke,Det ser ut på stormar och aldrig skakas;Det är stjärnan på varje vandrande bark,Vars värde är okänt, även om hans höjd tas.Älska oss inte Time dåre, men rosiga läppar och kinderInom hans böja skäran kompass komma;Kärlek förändrar inte med sina korta timmar och veckor,Men bär det ut ända till kanten av undergång.Om detta är fel och på mig visat,Jag har aldrig writen, eller ingen människa någonsin älskat.
		-- Walt Kelly

%
Låt oss gå då du och jagmedan natten läggs ut mot himlensom ett utstryk av senap på en gammal pork pie."Trevlig dikt Tom. Jag har idéer till förändringar men varför inte komma över?"
		-- Ezra

%
Låt oss gå genom vissa halv öde gator,De muttra retreatsAv oroliga nätter i en-natt billiga hotellOch sågspån restauranger ostronskal:Gator som följer som en mödosam argumentAv smygande intentAtt leda dig till en överväldigande fråga ...Åh, inte frågar, "Vad är det?"
		-- T. S. Eliot, "Love song of J. Alfred Prufrock"

%
Låt oss behandla män och kvinnor väl;Behandla dem som om de vore verkliga,Kanske de är.
		-- Ralph Waldo Emerson

%
Livet är som en burk sardiner.Vi är alla oss, letar efter nyckeln.
		-- Beyond the Fringe

%
Livet är vad som händer med dig när du upptagen med att göra andra planer.
		-- John Lennon, "Beautiful Boy"

%
Lyft varje röst och sjungaTill jord och himmel ring,Ring med harmonier av frihet;Låta vår glädje upphovHög som lyssnings himmel,Låt det ljuda högt som den rullande havet.Sjunga en sång full av tron ​​att det mörka förflutna har lärt oss.Sjunga en sång full av hopp om att den nuvarande har köpt oss.Vänd mot soluppgången i vår ny dag börjat,Låt oss marschera på till segern är vunnen.
		-- James Weldon Johnson

%
Lätta upp, medan du fortfarande kan,Inte ens försöka förstå,Bara hitta en plats för att göra din monter,Och ta det lugnt.
		-- The Eagles, "Take It Easy"

%
Som majs i ett område jag skära ner dig,Jag kastade den sista punch alldeles för hårt,Efter år av att gå stadigt, ja, jag tyckte det var dags,Att kasta i min hand för en ny uppsättning kort.Och jag kan inte ta dig att dansa ut på helgen,Jag tänkte att vi skulle målas alltför mycket i denna stad,Och jag försökte att inte titta när jag gick till min vagn,Och jag visste då jag hade förlorat vad som borde ha funnits,Jag visste då jag hade förlorat vad som borde ha funnits.Och jag känner mig som en kula i pistolen av Robert FordJag är så låg som en betald mördare ärDu vet att jag fryser som en hyrd svärd.Jag skäms vi inte kan lappa ihop det,Du vet att jag kan inte tänka klart längreDu gör mig känns som en kula, honung,en kula i pistolen av Robert Ford.
		-- Elton John "I Feel Like a Bullet"

%
"Linjer som är parallella träffas på Infinity!"Euclid flera gånger, hetsigt, manade.Tills han dog, och så nådde denna närhet:i det han fann att de förbannade saker gick isär.
		-- Piet Hein

%
Lisp, Lisp, Lisp Machine,Lisp Machine är kul.Lisp, Lisp, Lisp Machine,Kul för alla.
		-- Piet Hein

%
Little Fly,Din sommar spel Om tanken är livetMin tank handen och styrka och andas,Har brush'd bort. Och de villTanke är död,Är jag inteEn fluga som dig? Då är jagEller Är icke En lycklig flugaEn man som jag? Om jag borEller om jag dör.För jag dansarOch dricka och sjunga,Tills någon blinda sidanSkall borsta mina vingar.
		-- William Blake, "The Fly"

%
Lizzie Borden tog en yxa,Och försatt det djupt in i VAX;Har du inte avundas människor somGöra alla de saker ___ DU vill göra?
		-- William Blake, "The Fly"

%
Logiker har men dåligt definieradeSom rationella mänskligheten.Logik, säger de, tillhör människan,Men låt dem bevisa det om de kan.
		-- Oliver Goldsmith

%
Louie Louie, jag måste gåLouie Louie, jag måste gåFin liten flicka hon väntar på migMe fånga fartyget för över havetMe seglar fartyget ensam Tre nätter och dagar mig segla havetMig aldrig tänker mig göra det hem mig att tänka på flicka ständigt(Kör) På skeppet jag drömmer hon därJag luktar ros i håretMe se Jamaica månen ovan (kör, gitarrsolo)Det kommer inte att dröja länge, jag ser min kärlekJag tar henne i mina armar och sedanMig berätta att jag lämnar aldrig igen
		-- The real words to The Kingsmen's classic "Louie Louie"

%
Kärlek i ditt hjärta var inte där för att stanna.Kärlek är inte kärlek tills du ge bort.
		-- Oscar Hammerstein II

%
Kärlek, som snabbt tände i en mild hjärta,grep här för mässan formensom togs från mig-och vägen för det afficts mig fortfarande.Love, som frikänner ingen älskade en från att älska,grep mig så starkt med glädje i honom,att, som ni ser, det lämnar inte mig även nu.Kärleken tog oss till ett dödsfall.
		-- La Divina Commedia: Inferno V, vv. 100-06

%
Margaret, du sörjerÖver Goldengrove unleaving?Blad, som saker av människan,Du, med din nya tankarTa hand om, kan du?Ah! som hjärtat blir äldreDet kommer att komma till sådana sevärdheter kallareEfter hand, och inte heller skona en suckÄven världar wanwood leafmeal lögnOch ändå kommer du att gråta och vet varför.Nu spelar ingen roll, barn, namnetSorg är fjädrar är densamma:Det är fördärv mannen föddes för,Det är Margaret du sörja för.
		-- Gerard Manley Hopkins.

%
Meanehwael, baccat meaddehaele, monstaer lurccen;Fulle få alltför många drincce, hie luccen för fyht.[D] en Hreorfneorht [d] HWR, son Hrwaerow [p] heororthwl,AEsccen aewful jeork att steop outsyd.[P] hud! Bashe! Krasch! Beoom! [D] e Bigge gyeEallum hans bon brak, byt näsan offe;Wicced Godsylla waeld på hans asse.Monstaer moppe fleor wy [p] eallum män i haelle.Beowulf i bacceroome fonecall bemaccen Waes;Hearen sond av ruccus Saed "Hwaet [d] e helle?"Graben sheold Strang ond swich-blaed ScharpSond feorth att fyht [d] e grimlic fiende."Me" Godsylla Saed "mac [d] e minsemete."Heoro cwyc geten heold wi [p] faemed halv-nelsonOND Flyng honom lic frisbe bac att fen.Beowulf magen upp till meaddehaele bar,Saed, "Ne foe slagen mie faersom cUNG-fu."Eorderen Cocca-colha YCE-coeld [d] e reol [p] Yng.
		-- Not Chaucer, for certain

%
De flesta människor de tycker dagtid,"Orsakar de vilja se strålande solen.De är upp på morgonen,off och en gående tills de är alltför trött för att ha roligt.Men när solen går ner,och the bright lights skina, har min dagtid bara börjat.Nu finns det två sidor till denna stora värld,och en av dem är alltid natt.Om du kan ta hand om verksamheten i solen, baby,Jag antar att du kommer att bli bra.Do not come söker mig att låna ut en hand.Mina ögon bara inte kan stå ljuset.För att jag är en nattuggla honung, sova hela dagen lång.
		-- Carly Simon

%
Mamma damm för att göra mig gammal,Att svepa mina kläder, den svarta natt;Att åldras min röst, en gammal HÅGs kackel;Att bleka håret, ett skrik av skräck;En vindstöt till fläkt mitt hat;En blixt att blanda det väl -Nu börjar din magiska stava!
		-- Walter Disney, "Snow White"

%
Min analytiker sa att jag var rätt ut ur mitt huvud,Men jag sade, "Kära Doktor, jag tror att det är du istället.Eftersom jag har fått en sak som är unikt och nytt,För att bevisa det jag kommer att ha sista skratt på dig."Orsak stället för ett huvud - Jag har två.Och ni vet två huvuden är bättre än en.
		-- Walter Disney, "Snow White"

%
Min Bonnie såg i en gastank,Höjden på dess innehåll för att se!Hon tände en liten match för att hjälpa henne,Åh, ta tillbaka min Bonnie till mig.
		-- Walter Disney, "Snow White"

%
Min räknare är min herde, jag vill inteDet låter mig exakt tio signifikanta siffror,och det leder mig i grundpotens till 99 siffror.Det vederkvicker min kvadratrötter och vägleder mig längs stigar flytandedecimaler för tydlighetens skull.Ja, tho jag går genom dalen överraskning frågesporter,Fruktar jag intet prof, för min kalkylator är där för att glädja mig.Det bereder en stockbord för att trösta mig, det bereder enbåge synd för mig i närvaro av mina lärare.Det annoints min läxa med rätt lösningar, mina interpole äröver.Visst skall både precision och noggrannhet följa mig alla dagar av mittliv, och jag skall bo i huset av Texas Instruments för evigt.
		-- Walter Disney, "Snow White"

%
Min älskling fru var alltid dyster.Jag dränkte henne i en tunna rom,Och så såg till att hon skulle stannaI bättre sprit natt och dag.
		-- Walter Disney, "Snow White"

%
Min kärlek går förbi som en dag i juni,Och han gör inga vänner av sorg.Han kommer att trampa hans galopperande rigadoonI vägen eller morrows.Han kommer att leva sina dagar där solstrålarna börjarInte heller kunde storma eller vind utrota honom.Min egen kära kärlek, är han hela mitt hjärta -Och jag önskar somebody'd skjuta honom.
		-- Dorothy Parker, part 3

%
Min kärlek, han är galen, och min kärlek, är han flotta,Och en vild ung trä sak födde honom!Sätten är rättvist att hans roaming fötter,Och himlen är solbelyst för honom.Som kraftigt söt mitt hjärta verkar hanSom doften av akacia.Min egen kära kärlek, är han alla mina drömmar -Och jag önskar att han var i Asien.
		-- Dorothy Parker, part 2

%
My My, Hey HeyRock and roll är här för att stanna Kungen är borta men han inte glömtDet är bättre att bränna ut Detta är historien om en Johnny RottenÄn att blekna bort Det är bättre att bränna ut än det är att rostaMin min, hey hey Kungen är borta men han inte glömtDet är ur det blå och i den svarta Hey hey, my myDe ger dig detta, men du betalar för att Rock and roll kan aldrig döOch när du är borta kan du aldrig komma tillbaka Det finns mer i bildenNär du är ur det blå än med blotta ögatOch i den svarta"My My, Hey Hey (Out of the Blue), Rust Never Sleeps"
		-- Neil Young

%
"Mitt namn är Sue! Hur gör du ?! Nu ska du dö!"Tja, jag slog honom hårt rätt mellan ögonen,Och han gick ner, men till min förvåning,Kom upp med en kniv och skära av en bit av mitt öra.Så jag åkte en stol tvärs över tänderna,Och vi störtade genom väggarna och in i gatorna,Kickin 'och en-gougin' i leran och blodet och öl.Nu ska jag berätta för dig, jag har kämpat hårdare män,Men jag verkligen inte kan komma ihåg när:Han sparkade som en mula och han bet som en krokodil.Men jag hörde honom skratta och sedan hörde jag honom svära,Och han gick för sin pistol, men jag drog mitt första,Och han satt där lookin på mig, och jag såg honom le.Han sade: "Son, är den här världen grov,Och om en man som går att göra det han mĺste vara tuff,Och jag visste att jag inte skulle vara där för att hjälpa dig på vägen.Så jag ger dig det namnet och jag sa adjö,Och jag visste att du skulle behöva få svårt eller dö,Och det är det namnet som har hjälpt till att göra dig stark!
		-- Johnny Cash, "A Boy Named Sue"

%
Min egen kära kärlek, är han stark och fetOch han bryr sig inte vad som kommer efter.Hans ord ring söt som en fals av guld,Och hans ögon lyser med skratt.Han är jublande som en flagga unfurled -Åh, en flicka, hon inte glömma honom.Min egen kära kärlek, är han all min värld -Och jag önskar att jag hade aldrig träffat honom.
		-- Dorothy Parker, part 1

%
Min penna är på botten av en sida,Vilket är klar här historien slutar;'Tis att önska det hade förr gjort,Men berättelser på något sätt förlänga när börjat.
		-- Byron

%
Min själ är krossad, min ande ömJag tycker inte om mig längre,Jag anmärka, gräl, klagar, ripa,Jag funderar på smala husJag ryser vid tanken på mänJag är på grund av att bli kär igen.
		-- Dorothy Parker, "Enough Rope"

%
Natur att allt fast gränserna passar,Och klokt bromsas stolt man låtsas intelligens.Som på marken medan här vinster hav,I andra delar lämnar breda sandslätter;Således i själen medan minnet råder,Den fasta makt förståelse misslyckas;Där strålar av varm fantasi spel,Minnets mjuka siffror smälta bort.
		-- Alexander Pope (on runtime bounds checking?)

%
Nära Studio Jean CocteauPå Rue des Ecolesbodde en gammal manmed en blind hundVarje kväll jag skulle se honomstyra hund tillsammanstrottoaren, hållaett fast grepp på koppelså att hunden inte skullestöter på en förbipasserandeIbland hunden skulle slutaoch titta upp mot himlenNär gubbenmärke till mig att titta på hundenoch han sade, "Oh, ja,denna en vetnär månen är ute,han kan känna det på hans ansikte "
		-- Barry Gifford

%
Neuroser är röda,Melancholia blå.Jag är schizofren,	Vad är du?
		-- Barry Gifford

%
New York fick olika sätt;Bara inte låta dig vara.
		-- The Grateful Dead

%
New York-- som lång horisont kommer jagFlyin 'in från London till din dörrNew York-- Lookin ner på Central ParkDär de säger att du bör inte vandra after dark.New York.
		-- Simon and Garfunkle

%
Därefter på en pall, har vi en syn att göra dig dregla.Sju oskulder och en mule, hålla det svalt, håller det svalt.
		-- ELP, "Karn Evil 9" (1st Impression, Part 2)

%
Nio meg för sekreterarna rättvisa,Sju meg för hackare knappa,Fem meg för grads i rökiga lyor,Tre meg för systemkällan;En skiva att styra dem alla,En disk för att binda dem,En disk för att hålla filerOch i mörkret mala dem.
		-- ELP, "Karn Evil 9" (1st Impression, Part 2)

%
Niospårs band och sju-track bandOch band utan några spår;Stretch band och snarley bandOch band blandas upp på ställningar -Ta tag i bandetOch dra av remsan,Och då kommer du vara säkerBandenheten kommer att hoppa.
		-- Uncle Colonel's Cursory Rhymes

%
Ingen gillar oss.Jag vet inte varför.Vi kan inte vara perfekt, vi ger dem pengar,Men vem vet vi försöker. Men är de tacksamma?Men runt, nej, de är elak,Även våra gamla vänner sätta oss ner. Och de är hatiskt.Låt oss släppa den stora, De respekterar inte oss,Och se vad som händer. Så låt oss överraska demVi kommer att släppa den stora,Och pulverisera dem.Asiens trångt,Europa är för gammal,Afrika är alldeles för varmt, kommer vi att spara Australien.Och Kanadas för kallt. Vill inte skada någon kängurur.Och Sydamerika stal vårt namn vi kommer att bygga en All-American nöjenLåt oss släppa den stora, parkera there--Det blir ingen kvar att skylla oss. De fick Surfin ', också!bom! går London,Och Boom! Paree.Mer utrymme för dig, Oh, hur fredliga det ska vara!Och mer utrymme för mig, kommer vi ställa alla gratis!Och varje stad, du ska bära en japansk kimono, babe;Hela världen runt, Det blir italienska skor för mig!Kommer bara vara en annan amerikansk stad. Alla hatar oss hur som helst,Så, låt oss släppa den stora nu.Låt oss släppa den stora nu!
		-- Randy Newman, "Drop the Big One"

%
Ingen gris bör gå sky diving under monsunFör detta är egentligen inte normen.Men om ett fett svin försöka sväva som en galning,Än sen då? Alla fläsk i en storm.Ingen gris bör gå sky diving under monsun,Det är riskabelt nog när vädret är fint.Men att ha en gris sväva när monsun doth brusetKasta ännu fler faror för svin.
		-- Randy Newman, "Drop the Big One"

%
Ingen vanligt papper i löpande bana kan anse att fraktal Puff -Han växte så fort ingen plottning pack kunde krympa honom tillräckligt långt.Sammanställer och simuleringar växte så snabbt tamaOch bytte ut alla sina datautrymme när Puff sköt sin stack ram.(Avstå)Puff, blev han så snabbt, medan andra rörde sig som sniglarOch mini-Puffs skulle abborre sig på sin gigantiska svans.Alla student hackare älskade att fraktal PuffMen DCS inte gillar Puff, och till slut sa, "Nog!"(Avstå)Puff används mer resurser än DCS kunde avvara.Operatören dödade Puff jobb - han inte bry sig.En dysterhet föll på hackare; det verkade vara i slutet,Men Puff fångade undantag, och växte från noll igen!(Avstå)Avstå:Puff fraktal draken skriven i C,Och frolicked medan processer kopplas in stordator minne.Puff fraktal draken skriven i C,Och frolicked medan processer kopplas in stordator minne.
		-- Randy Newman, "Drop the Big One"

%
"Inget program är perfekt"De sa med en axelryckning."Kundens happy--Vad är en liten bugg? "Men han var fast besluten, sedan ändra två, sedan ytterligare tre,De andra gick hem. Som år följde år.Han grävde ut flödesschemat och främlingar skulle kommentera,Givna, ensam. "Är det killen fortfarande här?"Natten gick in i morgon. Han dog på konsolenRummet var rörigare av hunger och törstMed kärn soptippar, käll listor. Nästa dag han begravdes"Jag är nära", muttrade han. Sidan nedåt, nio kant först.Kedjan rökning, kallt kaffe, och hans fru genom tårarnaLogik, avdrag. Accepterat sitt öde."Jag har det!" ropade han, sade "Han är inte riktigt gått,"Bara ändra en instruktion." Han är bara arbetar sent. "
		-- The Perfect Programmer

%
Ingen sten så hårt men att en liten vågKan slå entré på tusen år.
		-- Tennyson

%
Knappt hade ogräs Allen PoeKom sin gamla Raven,då han började sin Old Crow.
		-- Tennyson

%
Nej, är hans sinne inte längre att hyraTill någon gud eller regering.Alltid hoppfull, men missnöje,Han vet förändringar är inte permanent -Men förändringarna är.
		-- Tennyson

%
Ingenting som är tvingade någonsin kan vara rätt,Om det inte kommer naturligt, lämna det.Det är vad hon sa när hon släckte ljuset,Och vi böjde ryggen som slavar i natten,Då sänkte hon sin vakt och visade mig ärrenHon fick från att försöka bekämpaSäger, åh, skulle du bättre tror det.[...]Väl ingenting som är verkligt är någonsin för gratisOch du behöver bara betala för det någon gång.Hon sagt det förut, sade hon till mig,Jag antar att hon trodde det fanns ingenting att se,Men samma gamla fyra imaginära väggarHon hade byggt för livin inneJag sade oh, du bara inte kan betyda det.[...]Väl ingenting som är tvingade någonsin kan vara rätt,Om det inte kommer naturligt, lämna det.Det är vad hon sa när hon släckte ljuset,Och hon kan ha varit fel, och hon kan ha varit rätt,Men jag vaknade med frost, och märkte att hon hade förloratSlöjan som täckte hennes ögon,Jag sade oh, du kan lämna den.
		-- Al Stewart, "If It Doesn't Come Naturally, Leave It"

%
Nu hat är den i särklass längsta nöje;Män älskar i all hast, men de avskyr på fritiden.
		-- George Gordon, Lord Byron, "Don Juan"

%
Nu lägger jag mig tillbaka till vila.Talarens tråkig; motivets djup.Om han skulle sluta innan jag vaknar,Ge mig en knuff för godhet skull.
		-- Anonymous

%
Nu lägger jag mig ner för att sovaJag ber den dubbla lås kommer att hålla;Maj ingen tegelsten genom fönstret paus,Och ingen råna mig tills jag vaknar.
		-- Anonymous

%
Nu lägger jag mig ner för att sova,Jag ber Herren min själ för att hålla,Om jag skulle dö innan jag vaknar,Jag kommer att gråta i vånda, "misstag !! misstag !!"
		-- Anonymous

%
Nu lägger jag mig ner för att studera,Jag ber Herren Jag kommer inte att gå nötaktig.Och om jag inte lära sig detta skräp,Jag ber Herren att jag inte kommer att kuggar.Men om jag gör, inte synd mig alls,Bara lägga mina ben i salen.Säg till min lärare jag har gjort mitt bästa,Sedan stapla mina böcker på mitt bröst.
		-- Anonymous

%
Nu är det dags att säga adjöTill alla våra företag ...M-I-C (se nästa vecka!)K-E-Y (Varför? Därför att vi gillar dig!)MUS.
		-- Anonymous

%
Nu låten börja! Låt oss sjunga tillsammansSol, stjärna, måne och dimma, regn och molnigt väder,Ljus på spirande blad, dagg på fjädern,Vinden på öppna backen, klockor på ljungen,Vassen vid skumma poolen, liljor på vattnet:Old Tom Bombadil och floden-dotter!
		-- J. R. R. Tolkien

%
Nu mina sextio år och tio,Tjugo kommer inte igen,Och ta från sjuttio fjädrar en poäng,Det lämnar mig bara femtio mer.Och eftersom att titta på saker i blomFemtio fjädrar är lite utrymme,Om skogen jag kommer att gåAtt se körsbär hängde med snö.
		-- A. E. Housman

%
Nu när dagen tröttnar mig,Min längtan önskanKommer att få mer vänligt,Som en trött barn, den stjärnklara natten.Händer, lämnar av dina handlingar,Märk väl, glömma alla tankar;Alla mina styrkorLängtar bara att sjunka in i sömnen.Och min själ, obevakat,Skulle skjuta i höjden på utbredda vingar,Att leva i natts magiska sfärDjupare, mer omväxlande.
		-- Hermann Hesse, "Going to Sleep"

%
Nu vad skulle de göra om jag seglade bara bort?Vem fan verkligen tvingade mig att lämna i dag?Runnin 'låg på berättelser om vad gjorde det en boll,Vad skulle de göra om jag gjorde inget landfall? "
		-- Jimmy Buffet, "Landfall"

%
Nu är det dags att ha några stora idéerNu är det dags att göra några bestämda beslutVi såg Buddha i en bar ner söderTalking politik och kärnklyvningVi ser honom och han är alla spolas upp -Går vidare in i kroppen av en skalbaggeSig redo för en lång lång krypaHan är inte ingenting - han är inte någonting alls ...Död och pengar gör sin poäng en gång merI form av Philosophical mördareMark och Danny ta bussen uptownDödliga änglar för verkligheten och passionHa mod här och nuInte ta något från halvfärdiga buddhasNär du tror att du fick det betalas i sin helhetDu har ingenting - du fick ingenting alls ...Vi är på väg och vi ute efter Buddha.Vi vet hans namn och han får inte komma undan.Vi är på väg och vi ute efter Buddha.Det skulle ta ett skott - att blåsa bort honom ...
		-- Shriekback, "Gunning for the Buddah"

%
O ge mig ett hem,Där buffeln strövar omkring,Där rådjur och antilop spela,Där sällan hörsEn nedslående ord,"Orsak Så kan en antilop säga?
		-- Shriekback, "Gunning for the Buddah"

%
O kärlek, kunde du och jag med ödet konspirerarFör att förstå detta tyvärr tingens ordning hela,Kan vi inte krossa det till bitarOch forma den närmare våra hjärtan önskan?
		-- Omar Khayyam, tr. FitzGerald

%
O smal som en pil-trollspö! O klarare än rent vatten!O vass av den levande poolen! Fair flod dotter!O fjäder tid och sommartid, och våren igen efter!O vinden på vattenfall, och löven "skratt!
		-- J. R. R. Tolkien

%
o! Vandrare i skuggad markförtvivlan inte! För att mörka de står,alla träslag finnas måste sluta äntligenoch se den öppna solen gå förbi:den nedgående solen, den uppgående solen,dagens slut, eller dagen börjat.För öst eller väst alla träslag måste misslyckas ...
		-- J. R. R. Tolkien

%
Observera yon plumed biped bra.För att aktivera sin captiva,Insättning på dess upphörande,En kvantitet av partiklar saltlösning.
		-- J. R. R. Tolkien

%
Av alla ord häxans undergångDet finns ingen så illa som vilka och vem.Mannen som dödar både som och vemKommer skrivas in i vår Vem är vem.
		-- Fletcher Knebel

%
Åh inte dagarna verkar lank och långNär allt går rätt och ingen går fel,Och är inte ditt liv extremt plattMed ingenting alls att klaga på!
		-- Fletcher Knebel

%
Oh ge mig din synd!Jag är på en kommitté Vi deltar och ändraVilket innebär att från morgon och brottas och försvaratill kväll, utan en slutsats i sikte.Vi ger och instämmer,Vi skjuta och demur, vi revidera agendanOch upprepa alla våra tankar. Med frekventa tilläggOch överväga en massa rapporter.Vi komponerar och föreslåVi antar och motsätter Men trots olika föreställningarOch punkterna förfarande är kul; Tas upp som motioner,Det är fruktansvärt lite blir gjort.Vi löser och befriar;Men vi aldrig lösa,Eftersom det är uteslutet för ossFör att få vårt utskottAtt sluta så här sång,Som stannar med en period, alltså.
		-- Leslie Lipson, "The Committee"

%
O Herre, vill du inte köpa mig en 4BSD?Mina vänner alla fick källor, så varför kan jag inte se?Kom du moby hackare, kom sjunga den med mig:Åt helvete med advokater från AT & T!
		-- Leslie Lipson, "The Committee"

%
"Åh," Melia, min kära, gör detta allt krona!Vem skulle ha trott jag skulle träffa dig i stan?Och varifrån detta verkliga plagg prosperi-ty? ""Åh, inte du vet att jag hade blivit förstört?" sade hon."Du lämnade oss i spillror, utan skor eller strumpor,Trött på att gräva potatis och Borrstart upp bryggor;Och nu har homosexuella armband och ljusa fjädrar tre! ""Ja: Det är hur vi klär när vi förstört", sade hon."Hemma i barton du sa 'dig' och 'du'Och `thik oon 'och` Theas oon' och 't'other; " men nuDu pratar ganska passar "ee för compa-ny!""En del polska vinns med en ruin", sade hon."Dina händer var som tassar sedan ditt ansikte blå och dysterMen nu är jag förhäxad av din känsliga kind,Och din lilla handskar passar som som på alla la-dy! ""Vi gör aldrig arbete när vi förstört", sade hon."Du brukade kalla hem-liv hag-ridit dröm,Och du skulle suck, och du skulle strumpa; men för närvarande du verkarAtt veta inte av glasvar eller melancho-ly! ""True. En är ganska livlig när förstört", sade hon."Jag önskar att jag hade fjädrar, en fin svepande klänning,Och en delikat ansikte, och kunde stötta om stan! ""Min kära - en rå land flicka, som du,Kan inte riktigt förväntar sig att. Du är inte förstört, "sade hon.
		-- Thomas Hardy

%
Åh, förresten, vilken Pink?
		-- Pink Floyd

%
Åh, ge mig ett hem,Där buffeln strövar omkring,Och jag ska visa dig ett hus med en riktigt rörig kök.
		-- Pink Floyd

%
Åh, ge mig ett ställe där gravitons fokusDär tre-body problem löses,Om mikrovågorna tona ner på tre grader K,Och förkylningsvirus aldrig utvecklats. (kör)Vi äter alger paj, vår vakuum är hög,Våra kullager är perfekt runda.Vår horisont är krökt, våra stridsspetsar är MIRVed,Och ett kilo väger ett halvt pund. (kör)Om vi ​​får slut på utrymme för vår spirande rasInga fler Lebensraum kvar för MenschNär vi är redo att börja, kan vi ta Mars isär,Om vi ​​bara hitta en tillräckligt stor skiftnyckel. (kör)Jag är trött på denna plats, det är bara McDonalds i rymden,Och leva upp här är ett hål.Säg till shiggies, "Do not cry", de kan kyssa mig farvälFör jag ska flytta nästa vecka till L4! (kör)KÖR: Home, hemma på LaGrange,Där rymdskrot alltid samlar in,Vi har, så det verkar, två av människans största drömmar:Solenergi och noll-gee sex.
		-- to Home on the Range

%
Åh, jag är en C programmerare och jag är okejJag muck med index och structs hela dagenOch när det fungerar, jag skrika hoo-rayÅh, jag är en C programmerare och jag är okej
		-- to Home on the Range

%
Åh, jag har halkat de sura band av jord,Och dansade himlen på skratt försilvrade vingarna;Sunward Jag har klättrat och anslöt sig till tumlande munterhetAv sol-split moln och gjort hundra sakerDu har inte drömt om -Grävmaskin och skjutit i höjden och svängdeHögt i den solbelysta tystnad.svävar därJag har jagat skrika vinden längs och kastadeMin ivriga hantverk genom fotlös salar luft.Upp, upp längs yrande, brännande blåJag har toppade vindpinade höjder med lätt nåd,Där aldrig lark, eller till och med örn flög;Och medan med tyst, lyft sinne Jag har beträddeDen höga untrespassed helighet utrymme,Sätt ut min hand och rörde vid Guds ansikte.
		-- John Gillespie Magee Jr., "High Flight"

%
Åh, är livet en härlig cykel av sång,Ett medley av extemporanea;Och kärlek är något som aldrig kan gå fel;Och jag är Marie av Rumänien.
		-- Dorothy Parker, "Comment"

%
Åh, hal Dee, kröp han ut ur havet.Han kan fånga alla de andra, men han kommer inte att fånga mig.Nej, han kommer inte att fånga mig, dumma ol 'slingrande Dee.Han kan fånga alla de andra, men AAAARRRRGGGGHHHH !!!!
		-- The Smothers Brothers

%
Åh, när jag var kär i dig,Då var jag ren och modig,Och miles runt undrar växteHur väl jag beter.Och nu fancy passerar,Och ingenting kommer att förbli,Och miles runt de kommer att säga att jagÄr ganska själv igen.
		-- A. E. Housman

%
Oh, ja, går livet vidare, långt efter det att spänningen i livin "är borta.
		-- John Cougar, "Jack and Diane"

%
Gamla mor Hubbard bodde i en sko,Hon hade så många barn,Hon visste inte vad jag ska göra.Hon flyttade till Atlanta.
		-- John Cougar, "Jack and Diane"

%
Gamla mor Hubbard gick till skåpetAtt hämta hennes dåliga dotter en klänning.När hon kom dit, skåpet var naknaOch så var hennes dotter, antar jag ...
		-- John Cougar, "Jack and Diane"

%
Old Tom Bombadil är en god kamrat,Klarblå kavajen är, och hans stövlar är gula.Ingen har någonsin fångat honom ännu, för Tom, är han mästare:Hans låtar är starkare låtar, och hans fötter är snabbare.
		-- J. R. R. Tolkien

%
På morgonen från en Bogart film, i ett land där de vände tillbaka tiden,Du går strosa genom folkmassan som Peter Lorre överväger ett brott.Hon kommer ut i solen i en sidenklänning kör som en akvarell i regnet.Bry dig inte om att be om förklaringar, kommer hon bara berätta att hon komI Year of the Cat.Hon ger inte tid för frågor, som hon låser upp armen i hennes,Och du följer "till din känsla av vilken riktning helt försvinner.Av de blå-kaklade väggar nära marknadsstånd finns en dold dörr hon    leder dig till.Dessa dagar, hon säger, jag känner mitt liv precis som en flod som rinner genomYear of the Cat.Jo, hon ser på dig så kallt,Och hennes ögon lysa som månen i havet.Hon kommer i rökelse och patchouli,Så du tar henne att hitta vad som väntar på insidanYear of the Cat.Tja, kommer morgon och du fortfarande med henne, men bussen och turister    är borta,Och du har kastat bort ditt val och förlorat din biljett, så du måste stanna på.Men trumma-beat stammar av natten kvar i takt med nyfödda dag.Du vet lite tid du är tvungen att lämna henne, men nu du ska boI Year of the Cat.
		-- Al Stewart, "Year of the Cat"

%
På det goda skeppet EnterpriseVarje vecka finns det en ny överraskningDär romulanerna lurarOch Klingonsen går ofta bärsärkagång.Ja, det goda skeppet EnterpriseDet finns spänning någonstans det flygerDär Tribbles spelarOch Nurse Chapel får aldrig sin väg.Se Kapten Kirk står på bryggan,Mr Spock är vid hans sida.Den veckovisa hot, ooh-oohDet blir stekt, spridda vitt och brett.Det är det goda skeppet EnterprisePå väg ut där faran liggerOch du bor i skräckOm du bär en skjorta som är röd.- Doris Robin och Karen Trimble The L.A. Filkharmonics,"The Good Ship Enterprise" till tonerna av "The Good Ship Lollipop"
		-- Al Stewart, "Year of the Cat"

%
Återigen fruktar gärning är gjort.Canon sover,hans allvetande öga skuggastill humant slump och omständighet.Fred råder på nytt o'er Pine Valley,men Canon sömn är oroliga.Akta, knappa dagar förbi Ides i juli.Otåliga händer vänta ivrigtatt förstå, att hållaknappa stunder av tidwrested från livet i den fullständigaära Canons makt;hålls fången av sin unblinking ögat.Tre gyllene klot stå vakt;en vardera till vägtullar i dag, timme, minuttills predestiny påbjuder hans reawakening.När det fruktade ögonblick arives,"Fråga inte för vem klockan klämtar,Det klämtar för dig. "Valley Pawn Shop idag "
		-- "I extended the loan on your Camera, at the Pine

%
Det var en liten nörd som älskade att läsa din e-post,Och sedan hämta tillbaka i-åtkomsttider för att få hackare av svansen,Och en gång när han avslutade läsning från sekreterarens spole,Han skrev en oförskämd avvisande till sin pojkvän (hur häftig!)Och detta som delivermail fungerade och han sprang sin backfstat,Han hörde ett fruktansvärt sprakande som råtta friterad i varmt fett,Och hårda fel förde ner systemet "därför han kan även skrika!Och bio bug'll ta din ner för EF du inte ser ut!Och när de var lite fling som skulle stryka genom uulog,Och när han gick till sin BLIT att natten för att spela på att vara Gud,OPS alla hörde honom ropa, och de till konsolen streckade,Men när de gjorde en ps -ut de hittade systemet kraschade!Åh, guiderna adb'd dumpar och gjorde systemet spår,Och arbetade i filsystemet 'til diskhuvudet var varm pasta,Men allt de någonsin hittats var detta: "panik: aldrig tvivel",Och bio bug'll krascha din box för EF du inte ser ut!När dagen är klar och månen kommer ut,Och du hör skrivaren gnälla och rk s verkar räkna,När den andra skrivbord är tomma och deras terminaler Glassy grå,Och lasten är bara 1,6 och du undrar om det ska bo,Du måste tänka filen skydd och inte snoka runt,Eller bio bug'll getcha och ta ner systemet!
		-- "I extended the loan on your Camera, at the Pine

%
En gång denna midnatt osammanhängande,Även om du funderade kännande och kristallin,Under många bruten och underordnadVolym av gnarly lore,Medan jag tjatade, nästan sång,Sudddenly kom en bilning,Som av någon ymnigt skulking,Skulking på min kammardörr.
		-- "I extended the loan on your Camera, at the Pine

%
En ljus söndag morgon, i skuggan av tornet,Genom Hjälp Office, jag sett mitt folk;När de stod där hungriga, jag stod där visslande,Detta land gjordes för dig och mig.Ingen levande någonsin kan stoppa mig,Som jag gå promenader denna frihet motorväg;Ingen levande någonsin kan göra mig att vända tillbaka,Detta land gjordes för dig och mig.Som jag gick promenader, såg jag en skylt där,Och på skylten det sa: "No Trespassing."Men å andra sidan, gjorde det inte säga någonting,Den sidan gjordes för dig och mig.[Om du någonsin undrat varför Arlo var så anti-establishment när hans pappaskrev sådana underbara patriotiska sånger, är svaret att du har intehört alla Woody låtar]
		-- Woody Guthrie, "This Land Is Your Land" (verses 4, 6, 7)

%
En dag,En galen meta-poet,Med inget att säga,Skrev en galen meta-diktDet började: "En dag,En galen meta-poet,Med inget att säga,Skrev en galen meta-diktDet började: "En dag,[...]sorts nära ".Var de ord som poeten,Slutligen valde,För att få sin galna dikt,Till någon form av nära ".Var de ord som poeten,Slutligen valde,För att få sin galna dikt,Till någon form av nära ".
		-- Woody Guthrie, "This Land Is Your Land" (verses 4, 6, 7)

%
En bra sak om musik,Tja, det hjälper dig att känna någon smärta.Så slog mig med musik;Hit mig med musik nu.
		-- Bob Marley, "Trenchtown Rock"

%
Ett piller gör dig större, och om du går jagar kaninerOch ett piller gör dig liten. Och du vet att du kommer att falla.Och de som mamma ger dig, Berätta dem en vattenpipa rökning larvInte göra något alls. Har gett dig samtalet.Fråga Alice Call AliceNär hon är tio fot lång. När hon var bara små.När män på schackbrädet när logik och proportionFå upp och berätta vart du ska gå. Fallit slarvig döda,Och du har bara haft någon form av och White Knight talarsvamp bakåtOch ditt sinne går låg. Och den röda drottningen förlorade huvudetFråga Alice Kom ihåg vad hasselmus sa:Jag tror att hon vet. Mata ditt huvud.						Mata ditt huvud.						Mata ditt huvud.
		-- Jefferson Airplane, "White Rabbit"

%
En anledning till varför George WashingtonHålls i en sådan vördnad:Han klandrade aldrig sina problemPå den tidigare administrationen.
		-- George O. Ludcke

%
En sak om det förflutna.Det är sannolikt att pågå.
		-- Ogden Nash

%
En toke över linjen, söta Mary,En toke över linjen,Sittin 'centrum i en järnvägsstation,En toke över linjen.Waitin 'för tåg som går hem,Hopin "att tåget är i tid,Sittin 'centrum i en järnvägsstation,En toke över linjen.
		-- Ogden Nash

%
Andra kvinnor cloyAptit de äter, men hon gör hungrigDär de flesta hon uppfyller.
		-- Antony and Cleopatra

%
Våra små system har sin dag,De har sin tid och upphöra att vara;De men trasiga lampor av dig.
		-- Tennyson

%
Våra fäder ålder var värre att våra grandsires ".Vi deras söner är mer värdelösa än de:så i vår tur ska vi ge världen en avkomma ännu mer korrupt.
		-- Quintus Horatius Flaccus (Horace)

%
Persiljaär gharsley.
		-- Ogden Nash

%
Payeen till en TwangderridaOre-Idapotatis.Om du vågade,Jag skulle be digatt gå grävaupp dina ides enligt brun-tubered himmel.där pitchforkeddu kommer att beDerrida?
		-- Ogden Nash

%
Plocka upp bitar av min söta krossade dröm,Jag undrar hur gamla människor är i kväll,Hennes namn var Ann och jag tusan om jag minns hennes ansikte,Hon lämnade mig inte veta vad man ska göra.Carefree Highway, låt mig glida iväg på dig,Carefree Highway, du sett bättre dagar,Morgonen efter blues, från mitt huvud ner till mina skor,Carefree Highway, låt mig glida iväg, glida bort, på dig ...Vrida tillbaka sidorna till de tider jag älskar bäst,Jag undrar om hon någonsin kommer att göra samma sak,Nu det som jag kallar livin 'är bara bein' nöjd,Med vetskap om jag fick ingen kvar att skylla.Carefree Highway, fick jag se dig, min gamla flamma ...Söka igenom fragment av min dröm krossades sömn,Jag undrar om de åren har stängt hennes sinne,Jag antar att det måste vara reslust eller tryin 'för att komma loss,Från den goda gamla trogna feelin 'vi en gång kände.
		-- Gordon Lightfoot, "Carefree Highway"

%
Rörsystem ned dalar vild,Piping låtar av trevliga glädje,På ett moln såg jag ett barn,Och han skrattar sade till mig:"Rör en sång om ett lamm!"Så jag leds med glatt mod."Piper, rör den låten igen;"Så jag leds Han grät höra.
		-- William Blake, "Songs of Innocence"

%
Plagiarize, plagiarize,Låt ingenmans arbete undvika ögonen,Kom ihåg varför goda Herren gjort dina ögon,Inte skugga dina ögon,Men plagierar, plagiarize, plagiera.Bara vara säker på att kalla det forskning.
		-- Tom Lehrer

%
Planet Claire har rosa hår.Alla träden är röda.Ingen dör någonsin där.Ingen har ett huvud ....
		-- Tom Lehrer

%
Vänligen stå för nationalsången:Australiensare allt, låt oss glädjas,För vi är unga och gratis.Vi har gyllene jord och välstånd för slitVårt hem är girt till sjöss.Vårt land är rikt på naturens gåvorAv skönhet rik och sällsynt.I historien sida, låt varje stegAdvance Australia Fair.I glada stammar låt oss sjunga,Advance Australia Fair.Tack. Du kan återuppta din plats.
		-- Tom Lehrer

%
Vänligen stå för nationalsången:Gud bevare vår Gracious Queen!Leve vår Noble Queen!God save the Queen!Skicka henne segrar,Glad och strålande,Lång tid att regera o'er oss!God save the Queen!Tack. Du kan återuppta din plats.
		-- Tom Lehrer

%
Vänligen stå för nationalsången:O CanadaVårt hem och hemlandSann patriot kärlekI alla dina söner kommandotMed glödande hjärtan ser vi dig stigaDen sanna norr stark och friFrån när och fjärran, O CanadaVi står på vakt för digGud hålla vårt land ärorika och gratisO Canada vi står på vakt för digO Canada vi står på vakt för digTack. Du kan återuppta din plats.
		-- Tom Lehrer

%
Vänligen stå för nationalsången:Åh, säger kan du se i gryningen tidiga ljusVad så stolt vi hyllades vid skymningen sista glimma?Vars breda ränder och ljusa stjärnor genom den farliga kampenO'er vallar vi såg var så galant streaming?Och raketerna "röda reflexer, bomberna spricker i luften,Gav bevis genom natten som vår flagga var fortfarande kvar.Åh, säg inte att stjärnspangled baner ännu vågO'er land of the free och hem för modiga?Tack. Du kan återuppta din plats.
		-- Tom Lehrer

%
Ström, som en förödande pest,Förorenar whate'er det berör ...
		-- Percy Bysshe Shelley

%
Trolig-Möjligt, min svarta höna,Hon lägger ägg i den relativa När.Hon inte lägga ägg i den positiva nuEftersom hon är oförmögen att postulera hur.
		-- Frederick Winsor

%
Föreslagna Country & Western låttitlarJag kan inte komma över dig, så jag utstyrseln och går runt till andra sidanOm du inte lämnar mig ensam, kommer jag hitta någon som kommerJag visste att du skulle begått en synd när du kom hem sent medDina strumpor utifrån och inJag är en kanin i strålkastarna på Your LoveInte sparka mina däck Om du inte är Gonna Take Me För en rittJag gillade dig bättre innan jag visste att du så braI Still Miss You, barn, men mitt mål är Getting BetterJag har röda ögon från dina White Lies och jag är blå hela tiden
		-- "Wordplay"

%
Föreslagna Country & Western låttitlarJag har inget emot om du ljuger för mig, så länge jag är inte Lyin AloneJag skulle inte ta dig till en Hundslagsmål Även om jag trodde du kan vinnaOm du lämnar mig, gå ut bakåt så jag tror att du är Comin 'InEftersom du lärt dig att Lip-Sync, jag är till ditt förfogandeVar min John Deere bryta ditt område, medan din Dear John Var	Krossar mitt hjärtaDo not Cry, Little Darlin ', Du Waterin "min ölTennis måste vara din racket, för kärlek betyder Nothin 'till digNär du säger att du älskar mig, du är full av katrinplommon, "Orsak LivingMed dig är PitsI Wanted din hand i äktenskap men allt jag fick var Finger
		-- "Wordplay"

%
Föreslagna Country & Western låttitlarHon är inte mycket att se, men hon ser bra ut genom botten av en GlassOm Fingeravtryck dök upp på hud, jag undrar vem är jag skulle hitta på digJag skäms över att vara här, men Inte skamset nog att lämnaDet är Commode Huggin 'Time In The ValleyOm du vill behålla öl Real kall, satte den bredvid min ex-frus hjärtaOm du får en känsla av att jag inte älskar dig, Känn igenJag skäms över att vara här, men inte skamset nog att lämnaDet är flaska mot Bibeln i kampen om pappas SoulMin fru sprang med min bästa vän, och jag säker saknar honomKlipp inte något mera Trä, baby, För jag ska är Comin 'Home med en lastJag älskade hennes ansikte, men jag lämnade henne bakom For You
		-- "Wordplay"

%
Annorlunda lösenord,Bomb ut, och försök igen.Försök att komma förbi inloggning,Vi hacking, dataintrång, hacking.Prova hans första fru flicknamn,Detta är mer än bara ett spel.Det är riktigt roligt, men precis samma,Det är hacking, dataintrång, hacking.
		-- To the tune of "Music, Music, Music?"

%
regnet faller där molnen kommasolen skiner där molnen gåmoln kommer bara och gå
		-- Florian Gutzwiller

%
Rakhyvlar smärta dig;Floder är fuktig.Syror fläcken dig,Och droger orsakar kramp.Vapen är inte tillåtet;Snaror ger.Gas luktar awful--Du kan lika gärna leva!
		-- Dorothy Parker, "Resume", 1926

%
Nå in tankar vänner,Och hitta de vet inte ditt namn.Pressa nallebjörn för hårt,Och titta fjädrarna spränga sömmarna.Tryck på blyinfattade med din kind,Och känna dess kyla på ditt blod.Hålla ett ljus till natten,Och se mörkret böja lågan.Riv masken av frid från Gud,Och höra bruset av själar i helvetet.Plocka en ros i kärlekens namn,Och titta på kronbladen curl och vissnar.Luta på den västra vinden,Och vet att du är ensam.
		-- Dru Mims

%
Reclaimer, skona trädet!Ta inte en enda bit!Den används för att peka på mig,Nu jag skydda den.Det var läsarens CONSSom gjorde det, parat med dot;Nu, GC, för nonce,Du skall återta det inte.
		-- Dru Mims

%
Kom ihåg att oavsett olycka kan vara din lott, kan det bara varasämre i Cleveland.
		-- National Lampoon, "Deteriorata"

%
Kom ihåg digAy, du dålig spöke medan minnet har en sitsI detta distraherad jordklotet. Kom ihåg dig!Ja, från bordet av mitt minneJag ska torka bort alla triviala förtjust poster,Alla sågar av böcker, alla former, alla tryck förbi,Att ungdomar och observation kopieras dit.
		-- William Shakespeare, "Hamlet"

%
Ta bort mig från detta land av slavar,Där alla är idioter, och alla är knaves,Där varje knekt och dåre är köpt,Ändå vänligt säljer sig för intet;
		-- Jonathan Swift

%
Roland var en krigare, från land midnattssolen,Med en Thompson pistol för uthyrning, kämpar för att göras.Affären gjordes i Danmark, på en mörk och stormig dag,Så han anges för Biafra, att ansluta sig till den blodiga striden.Genom sextiosex och sju, kämpade de Kongo krig,Med sina fingrar på sina triggers, knä djupt i gore.Dagar och nätter de kämpade, det Bantu på knä,De dödade tjäna sitt uppehälle, och att hjälpa den kongolesiska.Roland Thompson skytt ...Hans kamrater kämpade bredvid honom, Van Owen och resten,Men av alla Thompson artillerister, Roland var bäst.Så C.I.A beslutade de ville Roland döda,Det son-of-a-tik Van Owen, blåste av Roland huvud.Roland den huvudlösa Thompson skytt ...Roland sökte kontinenten, för mannen som hade gjort honom.Han fann honom i Mombasa, i en bar rum dricka gin,Roland syftar hans Thompson pistol, han sa inte ett ord,Men han blåste Van Owen kropp därifrån till Johannesburg.Den eviga Thompson skytt, fortfarande vandrar genom natten,Nu är det tio år senare, men han stillbilder håller upp kampen.I Irland, i Libanon, Palestina, i Berkeley,Patty Hearst ... hörde brast ... av Rolands Thompson pistol, och köpte den.
		-- Warren Zevon, "Roland the Headless Thompson Gunner"

%
Romeo var rastlös han var redo att döda,Han hoppade ut genom fönstret för att han inte kunde sitta stilla,Juliet väntade med ett skyddsnät,Sade "inte begrava mig för att jag är inte död ännu".
		-- Elvis Costello

%
Rosor är röda;Viol är blå.Jag är schizofren,Och så är jag
		-- Elvis Costello

%
Lördag natt i Toledo Ohio,Är som att vara någonstans alls,Under hela dagen hur timmar rusar förbi,Du sitter i parken och du tittar på gräset dör.
		-- John Denver, "Saturday Night in Toledo Ohio"

%
Säg det med blommor,Eller säg det med mink,Men vad du än gör,Säg det inte med bläck!
		-- Jimmie Durante

%
Säg många kameror fokuserade t'us,Våra medelålders skott gör oss rättvisa.Ingen rättvisa, snälla, förbannelse ye!Vi vill verkligen nåd:Du ser, 'tis rättvisa, äcklar oss.
		-- Thomas H. Hildebrandt

%
Säg min kärlek är enkelt haft,Säga att jag bitit rå med stolthet,Säga att jag är alltför ofta ledsen -Fortfarande se mig vid din sida.Säga att jag är varken modig eller ung,Säger jag uppvakta och dalta omsorg,Säg djävulen rörde min tunga -Du har fortfarande mitt hjärta att bära.Men säg mina verser inte skanna,Och jag får mig en annan man!
		-- Dorothy Parker, "Fighting Words"

%
Säga! Du har träffat en hög med trouble--Byst i affärer, förlorat din fru;Ingen bryr sig ett öre om dig,Du bryr dig inte ett öre för livet;Otur har hopp berövad dig,Hälsa misslyckas, önskar att du hade die--Varför du har fortfarande solen vänsterOch den stora blå himmel.
		-- R. W. Service

%
Science, Double Feature.Frank har byggt och förlorat sin varelse.Mörkret har erövrat Brad och Janet.Tjänarna gått till en avlägsen planet.Wo, oj, oj, oj.Vid sent på kvällen, dubbel funktion, bildspel.Jag vill gå, oj, oj, oj.Till sent på kvällen, dubbel funktion, bildspel.
		-- Rocky Horror Picture Show

%
Vetenskap! sant dotter till Old Time du konst!Som alterest allt med dina peering ögon.Varför preyest du alltså på poetens hjärta,Gam, vars vingar är tråkiga verkligheten?Hur skulle han älska dig? eller hur bedömer dig vis?Som wouldst inte lämna honom i hans vandrandeAtt söka efter skatt i juvel himmel,Även om han skjutit i höjden med en oförskräckt vinge?Har du inte dras Diana från sin bil?Och drivit Hamadryad från vedenAtt söka ett skydd i vissa lyckligare stjärna?Har du inte rivit Najaden från sin översvämning,Den Elfin från det gröna gräset, och från migDen sommardröm under tamarind trädet?
		-- Edgar Allen Poe, "Science, a Sonnet"

%
Scintillate, scintillate, metallkorn vivific,Fain hur jag pausar vid din natur specifik,Högdraget balanserande i etern rymlig,Mycket liknar en pärla kolhaltiga.Scintillate, scintillate, metallkorn vivific,Fain hur jag pausar vid din natur specifik.
		-- Edgar Allen Poe, "Science, a Sonnet"

%
Repa skivorna, dumpa kärnan stänga av den, dra ur kontaktenRulla banden över golvet, Ge kärnan en extra bogserbåtOch systemet kommer att krascha. Och systemet kommer att krascha.Teletypes krossas till bitar. Mem'ry kort, en och alla,Ge omfattningar några otäcka träffar kasta ut halvvägs ner i korridorenOch systemet kommer att krascha. Och systemet kommer att krascha.Och vi har också funnit Vänd bara en switchNär du slår på strömmen ned, och lamporna kommer att upphöra att ryckaDu vänder diskläsare i papperskorgen. Och bandenheter kommer att falla sönder						på ett ögonblick.Åh, det är så mycket roligt, när CPUNu processorn inte kommer att köra Kan skriva ut ingenting men "foo"Och systemet kommer att krascha. Systemet kommer att krascha.
		-- To the tune of "As the Caissons go Rolling Along"

%
Förförd, snarkade lurvig Samson.Hon scissored korta. Hårt klippt,Snart fjättrade slav, suckade Samson,Tyst intrigerande,Sightlessly sökerNågra vilde, spektakulära självmord.
		-- Stanislaw Lem, "Cyberiad"

%
Söka svärdet som var bruten:I Imladris bor den;Det skall råd tasStarkare än Morgul-stavar.Det ska visas en tokenDet Doom är nära till hands,För Isildurs Bane skall väckas,Och Halfling ut skall stå.
		-- J. R. R. Tolkien

%
Hon frågade mig, "Vad är ditt tecken?"Jag blinkade och svarade "Neon"Jag trodde jag skulle blåsa henne ...
		-- J. R. R. Tolkien

%
Hon förblindade mig med vetenskap!
		-- J. R. R. Tolkien

%
Hon kan döda alla dina filer;Hon kan frysa med rynkad panna.Och en våg av handen ger hela systemet ner.Och hon arbetar på sin kod till tio efter tre.Hon bor som en fladdermus, men hon är alltid en hacker för mig.
		-- Apologies to Billy Joel

%
Hon stod på spårenVinka armarnaLeder mig till det tredje järnvägs chockSnabb som en blinkningHon ändrade sigHon gav mig en nattDet är allt det varVad kommer det att ta tills jag slutarskojar självSlösar min tidDet finns inget annat jag kan göra"Orsak Jag gör allt för LeynaJag vill inte ha någon ny"Orsak Jag lever allt för LeynaDet finns ingenting i det för dig"Orsak Jag ger det till Leyna
		-- Billy Joel, "All for Leyna" (Glass Houses)

%
SHIFT TILL VÄNSTER!Förskjutning åt höger!POP UP trycka ner,BYTE, BYTE, BYTE!
		-- Billy Joel, "All for Leyna" (Glass Houses)

%
Flyttas till vänster,Flyttas till höger,Mask in, maskera,BYTE, BYTE, BYTE !!!
		-- Billy Joel, "All for Leyna" (Glass Houses)

%
Eftersom jag skada min pendelMitt liv är allt oberäkneligt.Min papegoja som var hjärtligNu sänder statisk.Mattan dog, kollapsade en palm,Katten håller gör bajs.Det enda som håller mig sanePratar med min sko.
		-- My Shoe

%
Sjunga hey! för badet vid slutet av dagenSom tvättar den trötta leran bort!En lommar är han som inte kommer att sjunga:o! Vatten Hot är en ädel sak!O! Sweet är ljudet av fallande regn,och bäcken som hoppar från backen till vanligt;men bättre än regn eller porlande bäckarär Water Hot som röker och ångar.o! Kallt vatten vi kan hälla på behovner en törstig hals och vara glad faktiskt;men bättre är öl, om dryck som vi saknar,och varma vattnet hälls ner på baksidan.O! Vatten är rättvist att hoppar på högi en fontän vitt under himlen;men aldrig gjorde fontän låter så sötsom stänker Varmvatten med mina fötter!
		-- J. R. R. Tolkien

%
Snövit! Snövit! O Lady klart!O drottning bortom den västra havet!O Lätt för oss att vandra härMitt i den värld av vävda träd!Gilthoniel! O Elbereth!Klart är dina ögon och ljust din andedräkt!	Snövit! Snövit! Vi sjunger till digI fjärran land bortom havet.O stjärnor som i Brun utan ÅrMed lysande hand av henne såddes,I blåsiga områden nu ljusa och klaraVi ser dig silver blomma blåst!O Elbereth! Gilthoniel!Vi minns fortfarande, vi som borI detta fjärran land under träden,Din starlight på västra Seas.
		-- J. R. R. Tolkien

%
Så mycketberorpåen rödhjulkärraglas medregnvattenbredvidden vitakycklingar.
		-- William Carlos Williams, "The Red Wheel Barrow"

%
Så, du bättre se upp!Du bättre inte gråta!Du bättre inte lyra!Jag säger dig varför,Jultomten kommer till byn.Han vet när du har sovit,Han vet när du är vaken.Han vet om du har varit dålig eller bra,Han har band till CIA.Så...
		-- William Carlos Williams, "The Red Wheel Barrow"

%
Så ... så du tror att du kan berättaHeaven från helvetet?Blå himmel från smärta? Har de få dig att handelnKan du berätta ett grönt fält Dina hjältar för spöken?Från en kall stålskena? Het aska för träd?Ett leende från en slöja? Varm luft för en sval bris?Tror du att du kan berätta? Klen tröst för förändring?Har du bytaEn promenad på en del i ett krigFör huvudrollen i en bur?
		-- Pink Floyd, "Wish You Were Here"

%
Soldater som vill vara en hjälteÄr praktiskt taget noll,Men de som vill vara civila,De kör in i miljoner.
		-- Pink Floyd, "Wish You Were Here"

%
Några av dem vill använda dig,Några av dem vill att användas av dig,... Alla letar efter något.
		-- Eurythmics

%
Några Primal termit knackade på trä.Och smakade det, och fann det bra.Och det är därför din kusin majFöll genom salongen golvet idag.
		-- Ogden Nash

%
Vissa säger att världen kommer att sluta i brand,Vissa säger i is.Från vad jag har ätit av lustJag håller med dem som förespråkar brand.Men om det skulle förgås två gånger,Jag tror jag vet nog av hatAtt säga att för destruktion, isÄr också braOch skulle räcka.
		-- Robert Frost, "Fire and Ice"

%
Ibland känner jag mig som jag blekna bort,Titta på mig, jag fick ingenting att säga.Gör inte mig arg med de saker spel som du spelar,Antingen tänds eller lämna mig ensam.
		-- Robert Frost, "Fire and Ice"

%
Ibland bor jag i landet,Och ibland jag bor i stan.Och ibland har jag en bra idé,Att hoppa i floden och drunkna.
		-- Robert Frost, "Fire and Ice"

%
Ibland ljusets alla skiner på mig,Andra gånger jag kan knappt se.På senare tid slår migVad en lång konstig resa det har varit.
		-- The Grateful Dead, "American Beauty"

%
Tala ungefär till din lilla pojke,Och slog honom när han nyser:Han bara gör det för att retaEftersom han vet att det retar.	Wow! Wow! Wow!Jag talar starkt för min pojke,Och slog honom när han nyser:För han kan verkligen njuta avPeppar när han vill!	Wow! Wow! Wow!
		-- Lewis Carrol, "Alice in Wonderland"

%
Tala ungefär till din lilla VAX,Och starta upp när den kraschar;Det vet att man inte kan slappna avEftersom personsökar thrashes!	Wow! Wow! Wow!Jag talar starkt till min VAX,Och starta upp när den kraschar;Trots alla mina favorit hackarMina jobb det alltid thrashes!	Wow! Wow! Wow!
		-- Lewis Carrol, "Alice in Wonderland"

%
På tal om Godzilla och annat som förmedlar skräck:Med en målmedveten grimas och en Mongo-liknande känslaHan kastar spinning hårddiskar i luften!Och han plockar upp en Vax och han kastar tillbakaNär han vadar genom labbet gör hemska ljud!Hjälplös användare med projekt på grundScream "Min Gud!" som han stomps på bandenheter, också!Å nej! Han säger Unix går för långsamt! Gå, gå, DECzilla!Oh, ja! Han kommer att ta upp VMS! Gå, gå, DECzilla! "* VMS är ett varumärke som tillhör Digital Equipment Corporation.* DECzilla är ett varumärke av ihåliga chokladharar av död, Inc.
		-- Curtis Jackson

%
Våren är här, Våren är här,Livet är käglor och livet är öl.
		-- Curtis Jackson

%
St Patrick var en gentlemansom genom strategi och stealthkörde alla ormarna från Irland.Här är en rost för hans hälsa -men inte alltför många toastingsså att du förlorar dig själv och sedanglömma den goda St Patrickoch se alla dessa ormar igen.
		-- Curtis Jackson

%
Stannade i sängen hela morgonen bara för att fördriva tiden,Det är något fel här, det kan inte vara mer förneka,En av oss förändras, eller kanske vi stannade bara försöker,Och det är för sent, baby, nu är det för sent,Även om vi verkligen har försökt att göra det,Något inuti har dött och jag kan inte dölja och jag kan bara inte fejka det ...Det brukade vara så lätt att leva här med dig,Du var lätta och luftiga och jag visste precis vad de ska göraNu kan du ser så olycklig och jag känner mig som en idiot.Det blir goda tider igen för mig och dig,Men vi kan inte bara hålla ihop, behöver du inte känna det också?Men jag är glad för vad vi hade och att jag en gång älskat dig ...Men det är för sent baby ...Det är för sent, nu älskling, det är för sent ...
		-- Carol King, "Tapestry"

%
Steg tillbaka, otrogna!Eller regnet aldrig kommer.Någon hålla elden brinnande, någon komma och slår på trumman.Du kanske tror jag är galen, du kanske tror att jag är galen,Men jag svär till dig, innan denna dag är slut,du folk är gonna se lite regn!
		-- Carol King, "Tapestry"

%
Konstiga saker görs för att vara nummer ettAtt sälja datorn Druiderna var företagare,IBM har deras strategem Och de byggde en granit lådaSom stadigt växer acuter, det spårade månen, varnade för monsuner,Och Honeywell konkurrerar som Hell, och prognos vårdagjämningenMen berättelsens felande länken Deras pris var rätt, deras framtidÄr systemet gammal Stonemenge säljs ljus,Av firman Druids, Inc. Prototypen säljs;Från Stonehenge webbplats sina bitar och byteSkulle fartyget för Celtic guld.De flyttfirma kom till lådan ramen;Den vägde en miljon ton!Trafiken folk tyckte det ett skämt Mannen talade sant, och därmed du(Vagnshjulen bara snurrade); En varning från tiderna;"De kommer ja sälja det" förmannen ditt lager kommer att glida om du inte kan levereraspottade, vad i din broschyr sidor."Bara lämna de vilda ogräs växer, se om det säljer utan klockorna"Det är Druid-typ, över utformade och strängar som ringer och darra;"Och magen upp de ska gå." Druid anseende gick ner i rännanEftersom de inte kunde leverera.
		-- Edward C. McManus, "The Computer at Stonehenge"

%
Lidande ensam existerar ingen som lider;Gärningen finns, men ingen görare därav;Nirvana är, men ingen söker det;Vägen finns, men ingen som reser den.
		-- "Buddhist Symbolism", Symbols and Values

%
Solen i natten, är alla tillsammans,Stigande i himlen, är liv för alltid.
		-- Brand X, "Moroccan Roll/Sun in the Night"

%
      / \ SUN av dem vill använda dig,     \\ \  / \ \\ / SUN av dem vill att användas av dig, / / \ / / // \ \ // \ \ // / SUN av dem vill att missbruka dig,  / / / \ /   / \\ \ SUN av dem vill att missbrukas ...     \ \\      \ /
		-- Eurythmics

%
Sweet sixteen är vackra Bess,Och hennes röst förändras - från "Nej" till "Ja".
		-- Eurythmics

%
System / 3! System / 3!Se hur det går! Se hur det går!Dess bildskärm förlorar så totalt!Den kör alla sina program i RPG!Den är gjord av vår favorit monopol!System / 3!
		-- Eurythmics

%
T: En stor monster, kallade han TROLL.Han vet inte rock, och han inte rullar;Dricka vin, och rök inga stogies.Han bara älskar att äta dem Roguies.
		-- The Roguelet's ABC

%
Ta en titt omkring dig, berätta vad du ser,En flicka som tror att hon är vanlig lookin hon har nyckeln.Om du kan få tillräckligt nära för att titta in i hennes ögonDet är något speciellt bakom bitterhet hon gömmer.Och du är rättvist spel,Man vet aldrig vad hon kommer att besluta, du är rättvist spel,Bara slappna av, njuta av åkturen.Hitta ett sätt att nå henne, gör dig själv en dåre,Men gör det med en liten klass, bortse från reglerna.För det här vet den nedersta raden, kunde inte få ett datum.Den fula ankungen slår tillbaka, och hon kommer att avgöra hennes öde.(Kör)De som du aldrig märker är de som du måste titta på.Hon är trevlig och hon är vänlig medan hon tittar på din grenen.Prova på samtal, är skvaller en lögn,Och att det finns tillräckligt hon tar dig hem och göra dig vill dö.(Kör)
		-- Crosby, Stills, Nash, "Fair Game"

%
Ta hjärta mitt i allt djupare dysterhet att din hund äntligen fåtillräckligt ost.
		-- National Lampoon, "Deteriorata"

%
Tan mig gömma sig när jag är död, Fred,Tan mig gömma sig när jag är död.Så vi garvade hans skinn när han dog, Clyde,Det hänger där på skjulet.Alla tillsammans nu...Bind mig känguru ner, sport,Binda mig känguru ner.Bind mig känguru ner, sport,Binda mig känguru ner.
		-- National Lampoon, "Deteriorata"

%
Berätta varför stjärnorna gör sken,Berätta varför murgröna garn,Berätta varför himlen är så blå,Och jag kommer att berätta just varför jag älskar dig.Kärnfusion gör stjärnor att lysa,FOTOTROPISM gör murgröna surrRayleighspridning gör himlen så blå,Könshormoner är därför jag älskar dig.
		-- National Lampoon, "Deteriorata"

%
Säg mig, O Octopus, ber jag,Är dessa saker armar, eller är de ben?Jag förundras över dig, bläckfisk;Om jag var du, skulle jag kalla mig oss.
		-- Ogden Nash

%
Terence, är denna dumma saker:Du äter dina proviant tillräckligt snabbt;Det kan inte bli mycket fel, 'tis klart,Att se den kurs du dricker din öl.Men Åh, bra Herre, versen du gör,Det ger en chap magen-värken.Kon, den gamla kon, är hon död;Det sover väl den behornade huvudet:Vi fattiga pojkar, 'tis vår tur nuAtt höra sådana låtar som dödade kon.Ganska väns 'tis att rimDina vänner till döds innan deras tid.Deppa, melankoli galen:Kom, rör en låt att dansa till, lad.
		-- A. E. Housman

%
Den känslan kom drygt mig.
		-- Albert DeSalvo, the "Boston Strangler"

%
Dessa pengar samtal,Jag ska inte förneka,Jag hörde det en gång,Det sade "Good-bye.
		-- Richard Armour

%
Reklambyrån SongNär kundens hoppande galen,Sätta sin bild i annonsen.Om han fortfarande skulle visa refraktär,Lägg en bild av sin fabrik.
		-- Richard Armour

%
Den allommjuk dominera stöten,Den tocsin i själen - middagsklockan.
		-- Lord Byron

%
Banken ringde för att berätta att jag är övertrasserat,Vissa freaks bränner kors på min gräsmatta,Och jag * kan inte * tro * det, alla Cheetos är borta,Det är bara en av dessa dagar!
		-- Weird Al Yankovic, "One of Those Days"

%
Banken skickade vårt uttalande i morse,Den röda färgen var en syn av stor vördnad!Deras siffror och gruvan kan ha en balanserad,Men min fru var alltför snabb på oavgjort.
		-- Weird Al Yankovic, "One of Those Days"

%
Bird of Time har men en liten väg att flyga ...och fågeln är på vingen.
		-- Omar Khayyam

%
Pojken stod på den brinnande däck,Äta jordnötter från Peck.Hans far kallade honom, men han kunde inte gå,För han älskade dessa jordnötter så.
		-- Omar Khayyam

%
Kamelen har en enda puckel;Den dromedar två;Annars tvärtom.Jag är aldrig säker. Är du?
		-- Ogden Nash

%
Karbonylen är polariserad,Delta änden är plus.Nukleofilen kommer således attack,Kolet kärna.Dessutom gör en alkohol,Typer finns men tre.Det är en bindning, för att motsvara,Från C till lysande C.
		-- Prof. Frank Westheimer, to "America the Beautiful"

%
Den gemensamma skarv, eller toppskarv,Lägger ägg inuti en papperspåse;Anledningen, ser du, utan tvekan,Är att hålla blixten ut.Men vad dessa ouppmärksam fåglarHar misslyckats med att märka är att besättningarBjörnar kan komma med bullarOch stjäla väskor att hålla smulor.
		-- Prof. Frank Westheimer, to "America the Beautiful"

%
Skillnaden mellan oss är inte mycket långt,cruising för hamburgare i pappas nya bil.
		-- Prof. Frank Westheimer, to "America the Beautiful"

%
Ögon Texas är på dig,All livelong dag;Ögon Texas är på dig,Du kan inte komma undan;Tro inte att du kan fly demFrån natten 'til tidigt på morgonen;Ögon Texas är på er'Til Gabriel blåser hans horn.
		-- University of Texas' school song

%
Trädgården är i sorg;Regnet faller svalt bland blommorna.Sommar rysningar tystPå sin väg mot sitt slut.Gyllene blad efter bladFaller från höga akacia.Sommar leenden, förvånade, svaga,I detta döende dröm om en trädgård.Under en lång stund, men i rosorna,Hon kommer att dröja på, längtan efter fred,och långsamtStäng hennes trötta ögon.
		-- Hermann Hesse, "September"

%
Blickar över cocktailsDet verkade vara så söttInte verkar ganska så amorösÖver Strimlad Vete
		-- Hermann Hesse, "September"

%
Den goda (jag är övertygad om, för en)Är men dålig lämnar ogjort.När ditt rykte är gjortDu kan leva ett liv roligt.
		-- Wilhelm Busch

%
Det goda livet var så svårfångadeDet fick mig verkligen nerJag var tvungen att återfå viss tillförsiktSå jag fick i kamouflage
		-- Wilhelm Busch

%
Den goda tiden närmar sig,Säsongen är till hands.När glatt klick på två-base lickKommer att höras över hela landet.Frosten dröjer kvar på jorden, ochBudless är träden.Men den glada ring röst vårenBärs på vinden.
		-- Ode to Opening Day, "The Sporting News", 1886

%
Graven är en fin och privat plats,men ingen, tror jag, gör det anamma.
		-- Andrew Marvell

%
Hoppet som fjädrar evigtSprings just upp din bakom.
		-- Ian Drury, "This Is What We Find"

%
Junior Gud leder nu rullenI listan över himlens kamrater;Han sitter i huset av hög kontroll,Och han reglerar sfärerna.Ändå gör han undrar, tror du att,Om, till och med i gudar gudomliga,Den bästa och klokaste kanske inte är de somSom har vältrade sig en stund med svin?
		-- Robert W. Service

%
De damer män beundrar, jag har hört,Skulle ryser vid en ond ord.Deras ljus ger en enda ljus;De skulle hellre stanna hemma på kvällen.De behöver inte hålla sig vaken till tre,Inte heller läsa erotisk poesi.De sanktionera aldrig det orena,Inte heller känner igen en ouvertyr.De krympa från pulver och från målarfärg ...Hittills har jag haft några klagomål.
		-- Dorothy Parker

%
Bladen var lång, gräset var grönt,Hemlock-umbels höga och rättvisa,Och i gläntan en ljus sågsAv stjärnor i skuggan skimrande.Tenn 'uviel var dans därTill musik av ett rör oseddaOch mot bakgrund av stjärnor var i hennes hår,Och i hennes kläder glimrande.Det Beren kom från berg förkylningar,Och förlorade han vandrade i bladen,Och där Elven-floden rulladeHan gick ensam och sörjande.Han kikade mellan odört bladenOch såg i konstigt blommor av guldVid sin mantel och ärmarna,Och hennes hår som skugga efter.Förtrollning läkte hans trötta fötterAtt över kullar var dömda att ströva omkring;Och tillbaka han skyndade, stark och flotta,Och grep på månstrålar glittrande.Genom vävda skogen i ElvenhomeHon flydde lätt på dans fötter,Och lämnade honom ensam fortfarande att ströva omkringI den tysta skogen lyssna.
		-- J. R. R. Tolkien

%
Lamporna är på,men du är inte hemma;din viljaär inte din egen;Ditt hjärta svettningar,Dina tänder slipa;ännu en kyssoch du kommer att vara min ...Du tror att du är immun mot grejer(Oh Yeah!)Det är närmare sanningen att säga att du inte kan få nog;Du vet att du kommer att ställas inför det,Du är beroende av kärlek! "
		-- Robert Palmer

%
Den lilla staden som tiden glömde,Där alla kvinnor är starka,De män är snygg,Och barnen över genomsnittet.
		-- Prairie Home Companion

%
Herren och jag är i ett får-herde relation, och jag är ien position negativ behov.Han prostrerar mig i en grön-bälte betesområde.Han leder mig riktnings parallellt med icke-brusande vattenflytande.Han återvänder till original tillfredsställelse min psykologiska makeup.Han slår mig på ett positivt beteende format för maximalprestige Hans identitet.Det ska verkligen sägas att trots att jag görambulatorisk framsteg genom umbragious inter-hill dödlighet platsen, skräckförnimmelser kommer inte att inledas i mig, på grund av para-Etiska fenomen.Din pastorala gånghjälpmedel och quadrupic pickup enhet presentera migi en pleasurific humöret.Du designar och producerar en näring bärande möbel typ strukturinom ramen för icke-kooperativa element.Du agerar ut en huvudrelaterad folk ritual som använder vegetabiliskt extrakt.Min dryck redskap upplever en volym kris.Det är en pågående avdragsgill faktum att din interrelationsempathetical och icke-ventious kapacitet kommer att behålla mig som derasrikta fokus under hela min icke-död period, och jag kommer att hahyresgäst rättigheter i bostadsenhet Herren på en permanent öppendeltid.
		-- Prairie Home Companion

%
Skaparna kan göraoch användarna kan använda,men fixeringsmedel måste fastställamed men minimala ledtrådar
		-- Prairie Home Companion

%
Mannen hade hon var snäll och renOch tillräckligt bra för varje dag,Men åh, kära vänner, du skulle ha settDen som kom undan.
		-- Dorothy Parker, "The Fisherwoman"

%
Morgonsolen när det är i ditt ansikte visar verkligen din ålder,Men som inte bry mig ingen; i mina ögon du är allt.Jag vet att jag håller dig roade,Men jag känner att jag används.Åh, Maggie, jag önskar att jag hade aldrig sett ditt ansikte.Du tog mig hemifrån,Bara för att rädda dig från att vara ensam;Du stal mitt hjärta, och det är vad som verkligen gör ont.Jag antar att jag kunde samla mina böcker och gå vidare tillbaka till skolan,Eller stjäla min pappas kö och göra en levande ur spela pool,Eller hitta mig en rock 'n' roll band,Som behöver en hjälpande hand,Åh, Maggie Jag önskar att jag hade aldrig sett ditt ansikte.Du gjorde ett första klassens narr av mig,Men jag är så blind som en dåre kan vara.Du stal min själ, och det är en smärta jag kan göra utan.
		-- Rod Stewart, "Maggie May"

%
Den flyttningen fingrar skriver; och, efter att ha writen,Går vidare: eller alla de Piety eller WitSka locka tillbaka för att avbryta en halv Line,Inte heller alla dina tårar tvätta bort ett ord av det.
		-- Rod Stewart, "Maggie May"

%
Nettot av lagen sprids så bred,Ingen syndare från dess svep kan dölja.Dess maskor är så fin och stark,De tar i varje barn av fel.O underbara väv av mysterium!Stora fiskar ensam flykt från dig!
		-- James Jeffrey Roche

%
Natten går snabbt när du soverMen jag är ute shufflin "för något att äta...Frukost på Egg House,Liksom våffla på grill,Jag är brända runt kanterna,Men jag är öm i mitten.
		-- Adrian Belew

%
Den L lama, han är en prästDe två L lamadjur, han är ett odjurOch jag kommer att satsa min siden pyjamasDet finns inte någon tre L lllama.hans avdelning svarade på något som liknar en "tre L lllama."
		-- O. Nash, to which a fire chief replied that occasionally

%
The Pig, om jag inte misstar mig,Ger oss skinka och fläsk och bacon.Låt andra tror att hans hjärta är stor,Jag tror att det dumt av grisen.
		-- Ogden Nash

%
Diktaren vars dålighet räddade hans livDen viktigaste poeten i sextonhundratalet var GeorgeVissna. Alexander Pope kallade honom "usel Wither" och Dryden sade om sinvers att "om de rimmade och rattled hela var väl".I vår egen tid, "The Dictionary of National Biography" konstaterar att hansarbete "är främst anmärkningsvärt för sin massa, smidighet och planhet. Den vanligtvissaknar äkta litterär kvalitet och ofta sjunker in imbecill knittel ".Hög beröm, faktiskt, och det kan fresta dig att njuta av en typiskgivande strof: Det är hämtad från "Jag älskade en jänta" och handlar omhögre känslor.Hon skulle mig "Honey" samtal,Hon hade - O hon skulle kyssa mig också.Men nu tyvärr! Hon har lämnat migFalero, Lero, toa.Bland andra detaljer i hans älskarinna som han valde att förevigavar hennes klokt val av skor.Femmor passade hennes sko.År 1639 den store poetens liv i fara efter hans tillfångatagande avrojalisterna under det engelska inbördeskriget. När Sir John Denham, denRojalistiska poet, hört talas om Wither förestående utförande, gick han till kungen ochbad att hans liv skonas. När frågade hans skäl, svarade John,"Därför att så länge Wither levde, Denham inte skulle redovisas ivärsta poet i England. "
		-- Stephen Pile, "The Book of Heroic Failures"

%
Predikanten, politikern, läraren,Var och en av dem en gång en barn.Ett barn verkligen är en underbar varelse.Vill jag en? God Forbiddie!
		-- Ogden Nash

%
Kaninerna The CowHär är en vers om kaniner kon av nötkreatur likar;Det betyder inte nämna deras vanor. Ena änden är mu, den andra, mjölk.
		-- Ogden Nash

%
Regnet det raineth på baraOch även om det orättvisa fella,Men framför allt på precis, därför attDen orättvisa stjäl bara paraply.
		-- Lord Bowen

%
Noshörningen är en hemtrevlig odjur,För det mänskliga ögat är han inte en fest.Farväl, farväl, du gamla noshörning,Jag stirrar på något mindre prepoceros.
		-- Ogden Nash

%
Vägen går någonsin på och påNer från dörren där det började.Nu långt framåt Vägen har gått,Och jag måste följa, om jag kan,Sysslar det med ivriga fötter,Tills det går något större sättDär många vägar och ärenden möts.Och vart då? Jag kan inte säga.
		-- J. R. R. Tolkien

%
Leende Våren kommer i glädje,Och buttre Winter flugor bistert.Nu kristallklart är de fallande vatten,Och Bonnie blått är klart.Färska o'er bergen bryter vidare på morgonen,Den ev'ning förgyller haven s svälla:Alla varelser glädje i solen återvänder,Och jag gläds i min bonnie Bell.Blommiga våren leder solig sommardag,Den gula hösten pressar nära;Sedan i sin tur komma dyster vinter,Till leende Spring igen visas.Således säsonger dans, liv framåt,Gamla tid och natur deras förändringar berätta;Men aldrig varierar, fortfarande oföränderliga,Jag älskar min Bonnie Bell.
		-- Robert Burns, "My Bonnie Bell"

%
Soldaten kom knackar på Drottningens dörr.Han sade: "Jag är inte slåss för dig längre."Drottningen visste att hon hade sett hans ansikte någonstans innan,Och sakta hon lät honom inne.Han sade: "Jag ser dig nu, och du är så mycket ung,Men jag har sett fler strider förlorade än jag har strider vunnit,Och jag har denna intuition att det är allt för ditt nöje.Och nu kommer du berätta varför? "
		-- Suzanne Vega, "The Queen and The Soldier"

%
Ljudet av substantiv är mestadels obunden.I staden ett substantiv kan bära en klänning,eller längre ner, kan klä en clown.Ett substantiv som är ljudet skulle aldrig clown,men osunda substantiv hoppa upp och ner.Ljudet av ett substantiv kan distrub plogning,och sedan, min kära, du skulle sättas i pund.Men snälla låt inte att få ner dig,anseende din klänning är tal om staden.
		-- A. Nonnie Mouse

%
Gatan predikanten såg så förbrylladNär jag frågade honom varför han kläddMed fyrtio pounds av rubrikerHäftade mot bröstet.Men han förbannade mig när jag visade honomJag sa, "Inte ens kan du dölja.Du ser, du är precis som mig.Jag hoppas att du är nöjd. "
		-- Bob Dylan

%
Solen skiner på havet,Lysande med all sin kraft:Han gjorde sitt bästa för att göraVågorna smidig och ljus -Och det var mycket märkligt, eftersom det varMitt i natten.
		-- Lewis Carroll, "Through the Looking Glass"

%
Tanke Polisen är här. De har kommitAtt sätta dig under hjärtstillestånd.Och eftersom de drar dig genom dörrenDe säger att du har missade testet.
		-- Buggles, "Living in the Plastic Age"

%
Spänningen är här, men det kommer inte att vara längeDet är bäst att ha din kul innan den rör sig längs ...
		-- Buggles, "Living in the Plastic Age"

%
Problemet med en kattunge är attNär det växer upp, det är alltid en katt
		-- Ogden Nash.

%
Problemet med digÄr problemet med mig.Fick två bra ögonMen vi fortfarande inte ser.
		-- Robert Hunter, "Workingman's Dead"

%
Sanningen du talar har inget förflutet och ingen framtid.Det är, och det är allt den behöver vara.
		-- Robert Hunter, "Workingman's Dead"

%
Sköldpaddan livs twixt pläterade däckSom i praktiken dölja sin kön.Jag tror att det smart av sköldpaddanI en sådan fix vara så fertila.
		-- Ogden Nash

%
Vädret är här, jag önskar att du var vacker.Mina tankar är inte alltför tydligt, men inte springa iväg.Min flickvän är ett hål; mitt jobb är för plikttrogen.Hell ingen är perfekt, vill du spela?Jag känner tillsammans idag!
		-- Jimmy Buffet, "Coconut Telegraph"

%
Vinden doth smakar så bitter sweet,Liksom Jaspar vin och socker,Det måste ha blåst genom någons fötter,Liksom de Caspar Weinberger.
		-- P. Opus

%
Den wombat bor över haven,Bland de avlägsna Antipodes.Han kan finnas på nötter och bär,Eller sedan igen, på missionärer;Hans avlägsna habitat utesluterAvgörande kunskap om hans humör.Men jag skulle inte engagera wombatI någon form av dödlig strid.
		-- "The Wombat"

%
Den värsta amerikanska PoetJulia Moore, "Sweet Singer of Michigan" (1847-1920) var så dålig attMark Twain sa hennes första bok gav honom glädje i 20 år.Hennes vers främst sysslar med våldsam död - den stora brandenChicago och gula febern epidemi visade naturliga ämnen för sin penna.Om döden var genom drunkning, genom anfall eller skenande släde, denformel var densamma:Har du hört talas om den fruktansvärda ödeMr P. P. Bliss och hustru?Av deras död jag kommer att beröra,Och även andra förlorade sina liv(I) Ashbula Bridge katastrof,Där så många människor dog.Även om du började någorlunda frisk i en av Julias dikter,chanserna är att efter några strofer du skulle vara på botten av enflod eller träffas av blixten. En kritiker av dagen sade hon var "värre änen Gatling gun "och i en tunn volym räknat 21 döda och nio skadades.Otroligt, några tidningar var kritiska av hennes arbete, ävenvilket tyder på att den söta sångerskan var "semi-kompetenta". Hennes svar varrättfram: "De redaktörer som har talat i denna skandalösa sätt har gåttbortom förnuftet. "Hon tillade att" litterärt verk är mycket svårt att göra ".
		-- Stephen Pile, "The Book of Heroic Failures"

%
Värsta versraderTill att börja med kan vi utesluta James Grainger lovande linje:"Kom, musa, låt oss sjunga om råttor."Grainger (1721-1767) inte har modet av hans övertygelse och raderasdessa ord på att upptäcka att hans lyssnare upplöst i spontanskratt det ögonblick de lästes upp.Ingen sådan motvilja drabbade Adam Lindsay Gordon (1833-1870) som varinspirerad av föremålet för krig."Flash! Flash! Bang! Bang! Och vi brann bort,Och grå taket rodnade och ringde;	Blixt! blixt! och jag kände hans kula flåSpetsen på mitt öra. Blixt! smäll!"Däremot, Cheshire ost provocerade John Armstrong (1709-1779):"... Det som Cestria sänder, envisa pasta fast mjölk ..."Medan John Bidlake styrdes av en medkänsla för grönsaker:"Den late morot sover sin dag i sängen,Krymplingar ärta ensam som inte kan stå. "George Crabbe (1754-1832) skrev:"Och jag var ask'd och tillstånd att gåAtt söka firman Clutterbuck och Co "William Balmford undersökt möjligheterna att religiös vers:"Så 'tis med kristna, Nature vara svagÄven i den här världen, riskerar att läcka ut. "Och William Wordsworth visade att han kunde göra det om han verkligen försökt närbeskriver en damm:"Jag har mätt det från sida till sida;Tis tre fot lång och två fot bred. "
		-- Stephen Pile, "The Book of Heroic Failures"

%
Den unga damen hade en ovanlig lista,Kopplat delvis en strukturell svaghet.Hon sätter inga förutsättningar.
		-- Stephen Pile, "The Book of Heroic Failures"

%
De, uh, snötäckta berg är som riktigt kallt, va?Och, um, slätter sträcka ut som min moms gördel, va?Det finns lotsa öl och munkar för alla, va?Så den sista att vara fredlig och allt är en stor idiot,va?Så stänga yer ansikte upp och torka yer mucklucks vid elden, va?Och drömma om flickor med sina höga balkar på, va?De kan vara kallt, men det är okej! Öl är bättre på det sättet!va?Skönhet!
		-- A, like, Tribute to the Great White North, eh?

%
Så här är till staden Boston,Staden skrik och stön.Där Cabots kan inte se Kabotschniks,Och Lowells inte kommer att tala till Cohns.
		-- Franklin Pierce Adams

%
Det finns dåliga tider precis runt hörnet,Det finns mörka moln hurtling genom himlenOch det är inte bra gnällOm en silverkantFör vi vet av erfarenhet att de inte kommer att rulla av ...
		-- Noel Coward

%
Det finns platser som jag kommer ihågHela mitt liv även om vissa har förändrats.Några evigt inte bättreNågra har gått och en del kvarstår.Alla dessa platser hade sina stunderMed älskare och vänner jag minns fortfarande.Vissa är döda och några bor,I mitt liv har jag älskade dem alla.Men av alla dessa vänner och älskare,Det finns ingen jämförelse med dig,Alla dessa minnen förlorar sin innebördNär jag tänker på kärlek som något nytt.Även om jag vet att jag kommer aldrig att förlora tillgivenhetFör människor och saker som gick före,Jag vet att jag ofta stanna upp och tänka på demI mitt liv har jag kommer att älska dig mer.
		-- Lennon/McCartney, "In My Life", 1965

%
Det finns konstiga saker gjorda i midnattssolAv de män som restprodukt för guld;De arktiska spår har sina hemliga berättelserDet skulle göra blodet att isas;Norrsken har sett konstiga platser,Men queerest de någonsin sågVar det natt på marge av sjön LebargeJag kremerade Sam McGee.
		-- Robert W. Service

%
Det finns i vissa levande själarEn kvalitet av ensamhet outsäglig,Så bra det måste delasSom företag delas av mindre varelser.En sådan ensamhet är min; så vet vid det härSom i oändlighetDet finns en ensammare än du.
		-- Robert W. Service

%
Det finns ingen anledning att vänta.Tåget stannade kör år sedan.Alla tidtabeller, broschyrer,De ljusa färgade affischer full av lögner,Promise rider till ett avlägset landSom inte längre existerar.
		-- Robert W. Service

%
Det finns något i pang förändringsMer än hjärtat kan bära,Olycka minnas lycka.
		-- Euripides

%
Det var en gång en sjöman som såg genom ett glasOch spionerade en rättvis sjöjungfru med skalor på hennes ... ön.Där måsarna flög över sitt bo.Hon kammade det långa håret som hängde över henne ... axlar.Och fick henne att kittla och klia.Sjömannen ropade "Det är en vacker ... sjöjungfru.En Sittin ute på klipporna. "Besättningen kom en kör, alla gripa sina ... glasögon.Och trångt fyra djup till järnväg.Alla ivriga att dela i denna fina del av ... nyheter...."Kasta ut en linje och vi ska lasso henne ... simfötter.Och snart vi kommer säkert att hittaOm sjöjungfrur är bättre före eller vara ... modigMina kära kamrater "Kaptenen ropade.Och förbanna med mjälte.Den här låten kan vara tråkigt, men det är absolut ren.
		-- Oscar Brand, "A Clean Song"

%
Det var en liten flickaSom hade en liten curlRätt i mitten av pannan.När hon var bra, hon var mycket, mycket braOch när hon var dåligt, var hon mycket, mycket populärt.
		-- Max Miller, "The Max Miller Blue Book"

%
Det finns en lärdom som jag måste komma ihågNär allt faller sönderI livet, precis som i kärleksfullDet finns en sådan sak som att försöka hårtDu mĺste sjungaSom du inte behöver pengarnaÄlska som du aldrig bli såradDu har gotta danceSom ingen tittarDet är gotta komma från hjärtatOm du vill att det ska fungera.
		-- Kathy Mattea

%
Det finns en spännande i beredskap för alla för vi är på väg att toastDet bolag som vi representerar.Vi är här för att muntra varje pionjär och även stolt skryta,Av detta man män vårt gedigna presidentNamnet T. J. Watson innebärEn mod ingen kan hejdaOch vi känner mig hedrad att vara här för att rosta IBM.
		-- Ever Onward, from the 1940 IBM Songbook

%
Det finns amnesi i en hangknot,Och komfort i yxan,Men det enkla sättet gift kommer att göra dina nerver slappna av.Det finns surcease i ett skott,Och sömn som kommer från ställningar,Men en praktisk utkast gift undviker hårdaste skatt.Du hittar vila på den heta knäböj,Eller gas kan ge dig pax,Men det närmaste hörnet kemisten har fred i paketerade staplar.Det finns tillflykt i kyrkan mycketNär du tröttnar på inför fakta,Och den jämnaste vägen är gift föreskrivs i vänligt quacks.Chorus: Med en * ugh * och en suck, och en kick av hälarna,Döden kommer tyst, eller det kommer med skriker -Men mest trivsamma platsen att hitta din slutÄr en kopp jubel från handen av en vän.
		-- Jubal Harshaw, "One For The Road"

%
Det finns lite att ta eller ge,Det finns lite i vatten eller vin:Denna levande, denna levande, denna levande,Var aldrig ett projekt av mina.Åh, är hårt kamp, ​​och gles ärFörstärkningen hos en vid toppen,För konst är en form av katharsis,Och kärlek är en permanent flopp,Och arbetet är provinsen nötkreatur,Och resten är för en mussla i ett skal,Så jag funderar på att kasta slaget -Vill du vänligen rikta mig till helvetet?
		-- Dorothy Parker

%
De sa att du hade visat det när de upptäckte våra resultatUngefär en månad innan. Deras hår började krypaBeviset var giltigt, mer eller mindre i stället för att förstå detMen något mindre än mer. Vi skulle köra sak genom PRL.Han sände dem ord som vi skulle försöka Do not tell en själ om allt dettaAtt passera där de hade misslyckats För det någonsin måste varaOch när vi har gjort, till dem En hemlig, hålls från alla andraDen nya bevis skulle skickas. Mellan dig och mig.Min uppfattning var att börja igenIgnorera alla hade de gjortVi vände det snabbt till kodFör att se om det skulle gå.
		-- Dorothy Parker

%
De gick rusar ner den motorväg,Trasslat runt och försvann.De brydde sig inte ... de var bara att dö för att få bort,Och det var liv i omkörningsfilen.
		-- Eagles, "Life in the Fast Lane"

%
De skulle inte lyssna på det faktum att jag var ett geni,Mannen sa "Vi fick alla som vi kan använda",Så jag har de stadigt-depressin "låg ner, mind-messin,Arbetar-på-biltvätt blues.
		-- Jim Croce

%
Thinks't du existens doth beror på tid?Det doth; men åtgärder är våra epoker; minaHar gjort mina dagar och nätter gängliga,Oändliga, och alla lika, som sand på stranden,Otaliga atomer; och en öken,Barren och kallt, på vilken de vilda vågorna bryter,Men ingenting vilar, spara slaktkroppar och vrak,Stenar, och saltsurf ogräs av bitterhet.
		-- Jim Croce

%
"Trettio dagar hath Septober,April, juni, och inte undra på.alla övriga har jordnötssmörutom min far som bär röda hängslen. "
		-- Jim Croce

%
Trettio vita hästar på en röd backe,Först de champ,Sedan stämpla,Då står de stilla.
		-- Tolkien

%
Denna ae nighte, detta ae nighte,Everye nighte och alle,Eld och slask och candlelyte,Och Christe motta thy Saule.
		-- The Lykewake Dirge

%
Detta här är flätverk,Emblem av vårt land.Du kan hålla den i en flaska;Du kan hålla den i handen.amen!
		-- Monty Python

%
Detta är för alla misshandlat assistenterOfödda och unbegot,För dem att läsa när de är i trubbelOch jag är inte.
		-- A. E. Housman

%
Detta är historien om bietVars kön är mycket svårt att seDu kan inte tala om han från honMen hon kan berätta, och så kan hanDen lilla biet är aldrig stillaHon har inte tid att ta p-pillerOch det är därför, i tider som dessaDet finns så många söner av bin.
		-- A. E. Housman

%
Detta är hur världen slutar,Detta är hur världen slutar,Detta är hur världen slutar,Inte med en smäll utan med ett kvidande.
		-- T. S. Eliot, "The Hollow Men"

%
Detta land är mitt land, och bara mitt land,Jag har ett hagelgevär, och du har inte fått en,Om du inte får ut, kommer jag blåsa huvudet av,Detta land är privat egendom.
		-- Apologies to Woody Guthrie

%
Denna sak allt slukar:Fåglar, djur, träd, blommor;Gnager järn, biter stål;Slipar hårda stenar till måltid;Dräper kung, fördärvar stad,Och slår högt berg ner.
		-- Apologies to Woody Guthrie

%
De som svettas i helvetets lågor, gå i ax blytunga, några trodde att deras inälvorHär är anledningen till att de föll: Lispeth fram sweetest vokaler.Även på jorden de bad i SAS, de erbjöd Dessa upp i berömPL / 1, eller annan råa, tänka allt detta stinkande hazeVulgar tunga. En Rapsody sung.Några Herren gjorde i högsta grad försöka Jabber av mindless hordenMontering alla sina grunder hex. Uppföljaren nästa gjorde håna herreTal som trätte som djävulens crable late uppföljare så enfangledHex som anges på Tower Babel Dess talarens läppar blev intrassladDen högsta steget. I sin propp.Eftersom i livet de bad så sjukOch erbjöd gud så snuskig matavfallNu svettas i helvetets lågorSvett från brist på APLSvett dynga!
		-- Apologies to Woody Guthrie

%
Även om jag respekterar att en hel delJag skulle få sparken om det var mitt jobbEfter att ha dödat Jason av ochOtaliga skrikande argonautsBlåsångare av vänlighetSom skyddsänglar detalltid näraBlå kanariefågel i utloppet av strömbrytareVem vakar över digGör en liten fågelholk i din själInte lägga alltför fin en punkt på denSäga att jag är den enda biet i din motorhuvGör en liten fågelholk i din själ
		-- "Birdhouse in your Soul", They Might Be Giants

%
Tre ringar för Elven-kings under bar himmel,Sju för dvärg-herrar i sina salar sten,Nio för Mortal Män dömda att dö,En för Dark Lord på hans mörka tronI delstaten Mordor där skuggor ligger.En ring att härska över dem alla, en ring för att hitta dem,En ring att föra dem alla och i mörkret binda demI delstaten Mordor där skuggor ligger.
		-- J. R. R. Tolkien, "The Lord of the Rings"

%
Kasta bort dokumentation och manualer,och användarna kommer att vara hundra gånger lyckligare.Kasta bort privilegier och kvoter,och användarna kommer att göra det rätta.Kasta bort egna och anläggningslicenser,och det kommer inte att finnas någon piratkopiering.Om dessa tre är inte tillräckligt,bara bo på din hemkatalogoch låt alla processer ha sin gång.
		-- J. R. R. Tolkien, "The Lord of the Rings"

%
Tickar ögonblicken som utgör en tråkig dagSlarva och avfall timmar på ett märkligt sättSparkar runt på en bit mark i din hemstadVäntar på någon eller något att visa dig vägenTrött på liggande i solen och sedan en dag hittar duStanna hemma för att titta på regnet tio år har fått bakom digDu är ung och livet är lång Ingen berättade när du ska köraOch det är dags att döda idag Du missade startskottetOch du kör och du kör för att komma ikapp med solen, men det sjunkerOch racing runt för att komma upp bakom dig igenSolen är densamma i ett relativt sätt men du är äldreKortare andetag och en dag närmare dödenVarje år blir kortare hänger på i tyst desperationär den engelska vägenaldrig tycks hitta tid Tiden är borta, är låten överPlaner som antingen kommit på skam trodde att jag skulle något mer att säga ...Eller en halv sida av klottrade linjer
		-- Pink Floyd, "Time"

%
Tiger fick jaga,Bird fick flyga;Man fick sitta och undra: "Varför, varför, varför?"Tiger fick sova,Fågel fick mark;Man fick berätta själv han förstå.
		-- The Books of Bokonon

%
Tim och jag en jakt gickVi hittade tre tärnor i ett tält,När de var tre, och vi var två,Jag bucked en och Timbuktu.
		-- the only known poem using the word "Timbuktu"

%
Tiden går, säger du?Ah nej!Tid kvar, * vi * gå.
		-- Austin Dobson

%
Tids tvättar renKärlek sår osedda.Det är vad någon sa till mig;Men jag vet inte vad det betyder.
		-- Linda Ronstadt, "Long Long Time"

%
'Tis drömmen om varje programmerare,Innan hans liv är gjort,Att skriva tre rader av APL,Och göra jävla saker och ting fungerar.
		-- Linda Ronstadt, "Long Long Time"

%
Till en snabb Young FoxVarför jogga utsökt bulk, fond galen vamp,Daft buxom jonquil, zephyr s gawky vice?Killen matas av arbete, quiz Joves xanthic lamp--Zow! Betänkligheter av deja vu gyp räv-kin tre gånger.
		-- Lazy Dog

%
att vara ingen annan än dig själv i en världsom gör sitt bästa dag och nattatt du som alla andrainnebär att bekämpa den svåraste stridennågon människa kan slåss ochaldrig sluta kämpa.
		-- e.e. cummings

%
Att koda det omöjliga kod, är detta min strävan -För att få upp en jungfru maskin, för att felsöka koden,Pop av ändlösa rekursion, oavsett hur hopplöst,Att grok vad som visas på skärmen, oavsett belastning,Att skriva dessa rutinerTill höger den unrightable bugg, utan tvekan eller paus,Oändligt rulla och thrash, att vara villiga att hacka FORTRAN IVAtt montera unmountable magtape, för en himmelsk orsak.För att stoppa den ostoppbara krasch! Och jag vet inte om jag bara ska vara santTill denna ärorika strävan,Och kön kommer att bli bättre för detta, det min kod körs CUSPy och lugn,Att en man, hånad och när det sätts på prov.bestämd att förlora,Fortfarande tvistade med hans sista tilldelningAtt skrota unscrappable kludge!
		-- To "The Impossible Dream", from Man of La Mancha

%
Att fela är mänskligt,Spinna kattdjur.
		-- Robert Byrne

%
Att fela är mänskligt, att spinna kattdjur.Att fela är mänskligt, två curs hund.Att fela är mänskligt, att moo nötkreatur.
		-- Robert Byrne

%
Allt finns det en säsong, en tid för varje pupose under himlen:En tid att födas, och en tid att dö;En tid att plantera och en tid att plocka vad planteras;En tid att döda, och en tid att läka;En tid att bryta ner, och en tid att bygga upp,En tid att gråta, och en tid att skratta;En tid att sörja och en tid att dansa;En tid att kasta bort stenar, och en tid att samla stenar;En tid att omfamna och en tid att avstå från att omfamna;En tid att vinna, och en tid att förlora;En tid att hålla och en tid att kasta bort;En tid att riva och en tid att sy;En tid att tiga och en tid att tala;En tid att älska, och en tid att hata;En tid av krig, och en tid av fred.Pred 3: 1-9
		-- Robert Byrne

%
Att stå och vara stilla,På Birkenhead borren,Är en förbannat tuff kula att tugga.
		-- Rudyard Kipling

%
Till vem morgonen är som nätter,Vad måste midnights vara!
		-- Emily Dickinson (on hacking?)

%
Att skriva en sonett måste du hänsynslöststrippar dina ord till nakna, villig kött.Då binder dem till en metafor eller tre,och ta med tvinga fram en tillfredsställande nät.Ordna dem din vilja, varje fot på plats.Du är befälhavaren här, och de slavarna.Nu piska dem att upprätthålla en konstant taktoch rytm som de står även i stavar.Ett ord som slår ingen glädje? Kasta ut!Vilken nytta är ord som driver inte till hjärtat?En lat frasen? Kassera den, skaka av tvivel,och välja mer foglig ord att ta sin del.En välutbildad sonett liv för att underhålla,genom samlag direkt till hjärnan.
		-- Emily Dickinson (on hacking?)

%
Tobak är en smutsig ogräs,Att från djävulen finns anledning;Det dränerar din plånbok, det bränner kläderna,Och gör en skorsten näsan.
		-- B. Waterhouse

%
Alltför häftigt att calypso,Alltför svårt att tango,För konstigt att Watusi
		-- The Only Ones

%
Troll satt ensam på sin plats av sten,Och mumsade och mumlade ett kalt gammalt ben;För många år hade han gnagt det nära,För kött var svårt att få tag på.	Gjord av! Gum av!I en grotta i bergen bodde han ensam,Och köttet var svårt att få tag på.Upp kom Tom med sina stora stövlar på.Sade han till Troll: "Be, vad youn?För det ser ut som shin O 'min nuncle Tim,Som bör vara en-lyin i kyrkogård.Caveyard! Paveyard!Detta många år har Tim varit borta,Och jag trodde att han var ljuger i kyrkogård. ""Min gosse", sade Troll, "detta ben jag stal.Men vad är ben som ligger i ett hål?Din nuncle var död som en klump o 'leda,Ovan Jag hittade hans skenbenet.Tinbone! Thinbone!Han kan avvara en aktie för en stackars trollFör han behöver inte hans skenbenet. "Sade Tom: "Jag kan inte se varför gillar o theeUtan axin "ledighet ska gå makin 'gratisMed skaftet eller smalbenet o 'min fars släkt;Så lämna den gamla ben över!Rover! Trover!Även döda han vara, det tillhör han;Så lämna den gamla bnone över! "
		-- J. R. R. Tolkien

%
Försök att inte.Do.Eller inte.Det finns inget försöka.
		-- J. R. R. Tolkien

%
"Twas bergen och eirie vägHar Mahwah i Patterson: "Akta sig Hopatcong, min son!Alla jersey var havet lundar, tänder som biter, naglarnaOch den röda banken Bayonne. att klo!Akta den bundna bäcken fågeln och skyHan tog sin belmar blad i hand: Kearney Communipaw ".Lång tid Folsom fiende han sökteTill vilade han med en bayway träd Och som i Nutley trodde han stod,Och stod en stund i tanken. Den Hopatcong med ögon flamma,Kom Whippany genom Englewood,Ett, två, ett, två, och genom Och Garfield som den kom.och genomDen belmar bladet gick Hackensack! "Och har du dödat Hopatcong?Han lämnade den döda och med det huvud Kom till mina armar, min Perth Amboy!Han gick Weehawken tillbaka. Hohokus dag! Soho! Rahway! "Han Caldwell i sin glädje.Har Mahwah i Patterson:Alla jersey var havet odlingarOch den röda banken Bayonne.
		-- Paul Kieffer

%
'Twas brillig och slithy TovesGjorde gyren och gimble i waben. "Akta sig Jabberwocken, min son!Alla mimsy var borogroves Käkarna som biter, klornaOch de Môme Raths outgrabe. att fånga!Akta Jubjub fågel,Han tog sin vorpal svärd i hand och sky frumious Bander! "Lång tid manxome fiende han sökte.Så vilade han av tumtum träd och som i uffish trodde stod hanOch stod en stund i tanken. The Jabberwock, med ögonen i brandKom whuffling genom Tulgey träEn! Två! En! Två! Och genom och och burbled som det kom!genomDen vorpal bladet gick snicker-mellanmål. "Hast du dödat Jabberwocken?Han lämnade den döda, och tog sitt huvud, kom till mina armar, min beamish pojke!Och gick galumphing tillbaka. Oh frabjous dag! Calooh! Callay! "Han chortled i sin glädje.'Twas brillig och slithy TovesGjorde gyren och gimble i waben.Alla mimsy var de borogrovesOch de Môme Raths outgrabe.
		-- Lewis Carroll, "Jabberwocky"

%
'Twas bullig och slithy mäklareKöpte och spela i vurm "Akta dig för Jabberstock, min son!Alla ljus var Dow Jones Stokers Kostnaden som biter, värdetGenom marknadens vrede unphased. som faller!Akta Econ'mist ord, och skyHan tog sin prognos svärdet i hand: Den falska Street o Walls "!Lång tid Boesk'some fiende han sökte -Sake likviditet, så d'intjänade han, och som i baisse trodde att han stodOch stod en stund i tanken. Den Jabberstock, med kläder av tweed,Kom waffling med sanningen för bra,Chip Black! Chip Blue! Och genom och yuppied bra med girighet!och genomPrognosen bladet gick snicker-mellanmål! "Och har du dödat Jabberstock?Det bet smutsen, och med sin skjorta, kom till min firma, V.P.ish pojke!Han gick studsade tillbaka. O stora pengar dag! Moolah! Bra spel! "Han köpte honom en Mercedes Toy.'Twas panik och slithy mäklareGjorde gyren och torktumlare i CrashAlla bräcklig var Dow Jones eldareOch mammon vrede dem bash!
		-- Peter Stucki, "Jabberstocky"

%
Twas FORTRAN som doloop gårGjorde logzerneg den ifthen blocketAlla kludgy var funktionen strömmarOch subrutiner adhoc.Akta runtime-bug min vänsqurooneg, den falska gotoAkta infiniteloopOch sky inprectoo.
		-- "OUTCONERR," to the scheme of "Jabberwocky"

%
'Twas midnatt på havet, Hennes barn var alla föräldralösa,Inte ett spårbundet var i sikte, Utom en en liten tot,Så jag klev in en cigarr butik som hade ett hem hela vägenAtt be dem om en ljus. Ovanför en ödetomt.Mannen bakom disken När jag såg genom ek dörrenVar en kvinna, gammal och grå, gick whale drifting av,Som används för att mixtra munkar Dess sex ben hängande i luften,På vägen till Mandalay. Jag kysste henne farväl.Hon sa "God morgon, främling", Denna berättelse en moralHennes ögon var torra med tårar, Som du tydligt kan se,När hon lade huvudet mellan fötterna Blanda inte din gin med whiskyOch stod så i år. På den djupa och mörka blå havet.
		-- Midnight On The Ocean

%
'Twas midnatt, och UNIX hackaGjorde gyren och gimble i deras grottaAlla mimsy var CS-VAXOch Cory Raths outgrabe."Akta programvaran röta, min son!Felen som biter, de jobb som thrash!Akta trasigt rör, och skyDen frumious systemet kraschar! "
		-- Midnight On The Ocean

%
'Twas natten innan krisen, och hela huset,Inte ett program arbetade inte ens en browse.Programmerarna var urvriden för mindless att bry sig,Veta chanser att cutover hade inte en bön.Användarna var inbäddat alla snug i sina sängar,Medan visioner av förfrågningar dansade i deras huvuden.När i lobbyn uppstod en sådan slammer,Jag sprang från min röret för att se vad som stod på.Och vad mina undrande ögon ska visas,Men en Super programmerare, omedveten att frukta.Snabbare än örnar hans program som de kom,Och han visslade och skrek och kallade dem vid namn;På uppdatering! På Lägg! På förfrågan! På bort!På batchjobb! På Utgående! På funktioner Complete!Hans ögon var glaserade över hans fingrar var mager,Från Helger och nätter framför en skärm.En blinkning i ögat och en vridning av huvudet,Snart gav mig att veta att jag hade inget att frukta ...
		-- "Twas the Night before Crisis"

%
'Twas natt segment av dygnsperiod   föregår den årliga Yuletide firandet, och   hela vår bostadsort,Kinetic aktivitet var inte i bevis bland   innehavare av denna potential, däribland   arter av inhemska gnagare kallas Mus musculus.Strumpor var minutiöst upphängd från den främre   kanten av den vedeldade caloric apparaten,I enlighet med vår föregripande nöje om en   hängande umgänget från en excentrisk   filantrop bland vars folkloric appelations   är den honorific titeln St. Nicklaus ...
		-- "Twas the Night before Crisis"

%
Tjugo två tusen dagar.Tjugo två tusen dagar.Det är inte mycket.Det är allt du har.Tjugo två tusen dagar.
		-- Moody Blues, "Twenty Two Thousand Days"

%
Två män såg ut från fängelsegaller,Man såg mud--De andra såg stjärnor.Låt mig få denna rätt: två fångar tittar ut genom fönstret.Medan en av dem var ute på alla leran - fick den andra en hiti huvudet.
		-- Moody Blues, "Twenty Two Thousand Days"

%
Tyger, tyger, brinnande ljus Där hammaren? Där kedjan?I skogarna i natten, i vilken ugn var din hjärna?Vad odödlig hand eller öga Vad städet? Vad fruktan greppVågar rama thy rädda symmetri? Våga sina dödliga skräck lås?Bränns i avlägsna djup eller himmel När stjärnorna kastade sina spjutDen grymma eld dina ögon? Och water'd himlen med sina tårarPå vilka vingar vågar han eftersträvar? Vågar han skrattar sitt arbete för att se?Vad handen vågar gripa branden? Vågar han som gjorde lammet göra dig?Och vad skuldra & vad konst Tyger, Tyger, brinnande ljusKan vrida senor av de hjärta? I skogarna i natten,Och när ditt hjärta började slå Vad odödlig hand eller ögatVad fruktan handen och vad rädsla fötter Våga rama din rädda symmetri?Kan hämta det från ugnen djupOch i dina hemska revben vågar brantI brunnen av sanguine ve?I vilken lera och i vilken mögelVar dina ögon raseri roll'd?
		-- William Blake, "The Tyger"

%
U: Det finns en U - en Unicorn!Kör rätt upp och gnugga dess horn.Titta på alla dessa punkter du förlorar!Umbra Hulks är så förvirrande.
		-- The Roguelet's ABC

%
Under den breda och tunga VAXGräv min grav och låt mig slappnaLänge har jag bott, och många mina hackaOch jag lägger mig ner med en vilja.Dessa är de ord som berättar hur:"Här ligger han som leds 64K,Fällde maskinen för nästan en dag,Och Rogue spelar en förfärlig stillastående. "
		-- The Roguelet's ABC

%
Under den breda och stjärnhimlen,Gräv min grav och låt mig ligga,Glad gjorde jag bor och gärna dö,Och lade mig ner med en vilja,Och detta vara versen som du grav för mig,Här ligger han där han längtade efter att vara,Home är sjömannen hem från havet,Och jägaren hem från berget.
		-- Robert Loius Stevenson, "Requiem"

%
Upp mot nätet, redneck mor,Mamma som har höjt din son så väl;Han är sjutton och Hackin "på en Macintosh,Flammande stavfel och russin "hell ...
		-- Robert Loius Stevenson, "Requiem"

%
Vid härden branden är röd,Under taket finns en säng;Men ännu inte trötta är våra fötter,Fortfarande runt hörnet vi kan mötaEn plötslig träd eller stående stenAtt ingen har sett men vi ensamma. Fortfarande runt hörnet kan det vänta  Träd och blommor och blad och gräs, en ny väg eller en hemlig port,  Låt dem passera! Låt dem passera! Och även om vi passera dem idag  Hill och vatten under himmel, morgon vi kan komma på detta sätt  Passera dem! Passera dem! Och ta de dolda vägar som körsMot månen eller solen,Home ligger bakom, världen framåt, Apple, tagg, och mutter och slån,Och det finns många vägar att beträda Låt dem gå! Låt dem gå!Genom skuggor till kanten av natten, sand och sten och pool och Dell,Fram till stjärnorna är alla lyser. Fare dig väl! Fare dig väl!Då värld bakom och hem framåt,Vi ska vandra tillbaka till hem och säng.  Mist och skymning, moln och skugga,  Bort skall blekna! Bort skall blekna!  Eld och lampa, och kött och bröd,  Och sedan till sängs! Och sedan till sängs!
		-- J. R. R. Tolkien

%
Tonlös det gråter,Vinglösa fladdrar,Otandade bett,Mouthless muttrar.
		-- J. R. R. Tolkien

%
Vulkan har en storhet som är dysterOch jordbävningar bara skrämma de dolts,Och för den som är vetenskapligtDet finns ingenting som är fantastisktI mönstret för en flygning av blixtar!
		-- W. S. Gilbert, "The Mikado"

%
Tuss någon makt giftie gie ossAtt se oursels som andra ser oss.
		-- R. Burns

%
Vakna nu mina glada grabbar! Vakna och höra mig ringer!Varm nu hjärta och lem! Den kalla stenen har fallit;Mörk dörren står bred; döda hand är bruten.Natten under natten flygs, och porten är öppen!
		-- J. R. R. Tolkien

%
Vakna upp alla ni medborgare, höra ert lands samtalInte till vapen och våld, men freden för alla och envar.Krossa ut hat och fördomar, rädsla och girighet och synd,Hjälp föra tillbaka sin värdighet, återställa sin tro igen.Arbeta hårt för en gemensam sak, låt inte vårt land falla.Gör henne stolt och stark igen, demokrati för alla.Ja, gör vårt land starkt igen, hålla vår flagga unfurled.Gör vårt land väl igen, respekteras av världen.Gör sin helhet och vacker, arbetar från sol till solen.Stå rak och arbets sida vid sida, eftersom det finns så mycket att göra.Ja, gör henne hela och vacker, förenade stark och fri,Vakna upp, alla ni medborgare, det är upp till dig och mig.
		-- Pansy Myers Schroeder

%
Vill berätta allt en berättelse 'bout en man vid namn Jed,En dålig bergsbestigare, höll knappt sin familj utfodras.Men så en dag han Shootin "någon mat,När upp genom marken kommit bubblin "rå - olja, är det;	svart guld; "Texas te" ...Väl nästa sak ya vet, gamla Jed en miljonär.Den fränder sade, "Jed flyttar därifrån!"De sa, "Californy är platsen ya oughta vara"Så de laddade upp lastbilen och de flyttade till Beverly - Hills, som är;Swimmin 'pooler; filmstjärnor.
		-- Pansy Myers Schroeder

%
Fanns det en tid då dansarna med sina fiolerI barns cirkusar kunde stanna sina bekymmer?Det fanns en tid kunde de gråta över böcker,Men tiden har satt sin maggot på deras spår.Enligt den båge av himlen de är osäkra.Vad har aldrig känt är säkrast i det här livet.Enligt skysigns de som inte har några armarHar renaste händer, och, såsom hjärtlösa spöketEnsam är oskadd, så den blinde mannen ser bäst.
		-- Dylan Thomas, "Was There A Time"

%
Tittar flickor går förbiDet är inte den senaste sakJag bara stod i en dörröppningJag försöker bara att göra någon meningAv dessa flickor som passerar genom en leende avlastar hjärtat som sörjerDe berättelser de berättar om män Kom ihåg vad jag saJag väntar inte på en dam jag inte väntar på en damJag bara väntar på en kompis jag bara väntar på en vän...Behöver inte en horaBehöver ingen spritBehöver inte oskuld präst Ooh, samlag och bryta hjärtanMen jag behöver någon jag kan gråta till Det är ett spel för ungdomarJag behöver någon att skydda Men jag väntar på en damJag bara väntar på en vänJag bara väntar på en vän
		-- Rolling Stones, "Waiting on a Friend"

%
Vi behöver inte ingen utbildning, vi behöver inte ingen tankekontroll.
		-- Pink Floyd

%
Vi behöver inte någon indirekthet Vi behöver ingen sammanställningVi behöver inte någon kontroll flödes Vi behöver ingen laststyrningInga data maskinskrivning eller deklarationer Ingen länk redigera för externa bindningarHallå! lämnade du listorna ensam? Hallå! lämnade du den källan ensam?Chorus: (Chorus)Oh Nej, det är bara en ren samtal LISP funktion.Vi behöver inte någon sida påverkande Vi behöver ingen tilldelningVi behöver inte ingen flödeskontroll Vi behöver inte några särskilda-noderInga globala variabler för utförande Ingen mörk bit-vändning för felsökningHallå! lämnade du args ensam? Hallå! lämnade du dessa bitar ensam?(Chorus) (Chorus)
		-- "Another Glitch in the Call", a la Pink Floyd

%
Vi måste komma ur denna plats,Om det är det sista vi någonsin gör.
		-- The Animals

%
vi kommer att uppfinna nya vaggvisor, nya låtar, nya handlingar av kärlek,Vi kommer att gråta över saker som vi brukade skratta &vår nya visdom kommer att föra tårar till ögonen av mildvarelser från andra planeter som var rädda för oss tills dess &i slutändan en sommar med vilda vindar &nya vänner blir.
		-- The Animals

%
Vi önskar dig en Hare KrishnaVi önskar dig en Hare KrishnaVi önskar dig en Hare KrishnaOch en Sun Myung Moon!
		-- Maxwell Smart

%
Vi är glada lilla Vegemites,Lika ljus som ljus kan vara.Vi alla njuta av vår VegemiteTill frukost, lunch och te.
		-- Maxwell Smart

%
Vi är Riddarna av runda bordetVi dansar whene'er vi kanVi gör rutiner och chorus scener Vi är riddare av det runda bordetMed fotarbete oklanderlig Våra föreställningar är formidabelVi äta bra här i Camelot Men många gångerVi äter skinka och sylt och Spam mycket. Vi har gett rimDet är ganska unsingableI krig vi tuff och kan, vi är opera galen i CamelotGanska outtröttlig Vi sjunger från membranet mycket.Mellan våra questsVi Paljett västarOch imitera Clark GableDet är ett upptaget liv i Camelot.Jag måste skjuta vagnen en hel del.
		-- Monty Python

%
Vi har provat varje snurrande utrymme moteOch räkna dess verkliga värde:Ta oss tillbaka till hemmen av mänPå den svala, gröna kullarna i jorden.Spännet sky ringerSpacemen tillbaka till sin handel.Alla händer! Står fast vid! Faller fritt!Och lamporna under oss blekna.Ut rida söner Terra,Långt driver dånande jet,Up hoppar loppet av Earthmen,Ut, långt, och framåt yet--Vi ber för en sista landningPå jorden som gav oss födelse;Låt oss vila ögonen på de ulliga himmelOch de svala, gröna kullarna i jorden.
		-- Robert A. Heinlein, 1941

%
Välkommen tillbaka, mina vänner, till showen som aldrig tar slut!Vi är så glad att du kunde närvara, komma in, komma in!Där bakom glaset finns en verklig grässtrå,Var försiktig när du passerar, röra sig längs, röra sig längs.Kom in, showen är på väg att starta,Garanterat att blåsa huvudet isär.Lugna, du får dina pengar är värt,Största show, i himlen, helvetet eller jord!Du måste se bildspelet! Det är en dynamo!Du måste se bildspelet! Det är rock 'n' roll!
		-- ELP, "Karn Evil 9" (1st Impression, Part 2)

%
Jo jag tittade på min klocka och det sade en 4:45,Rubriken skrek att jag fortfarande var vid liv,Jag kunde inte förstå det, jag trodde jag dog i går kväll.Jag drömde att jag hade varit i en gränsstad,I en liten cantina att pojkarna hade funnit,Jag var desperat att dansa, bara för att gräva den lokala ljud.När kom en senorita,Hon såg så bra att jag var tvungen att träffa henne,Jag var redo att närma sig henne med min engelska charm,När hennes mässing välvda pojkvän tog mig i armen,Och han sade, växer några funk egen, amigo,Odla någon funk egen.Vi har inte som att med gringo kampen,Men det kan finnas en död i Mexiko ikväll....Ta mitt råd, ta nästa flyg,Och växa lite funk, öka din funk hemma.
		-- Elton John, "Grow Some Funk of Your Own"

%
Tja, infall ger pengar till regeringen!Kunde lika gärna ha lagt ner i avloppet.Fancy ger pengar till regeringen!Ingen kommer att se saker igen.Jo, de har ingen aning om vad pengar är för -Tio till en de ska starta ett nytt krig.Jag har hört en hel del dumma saker, men Lor "!Fancy ger pengar till regeringen!
		-- A. P. Herbert

%
Tja, jag vet inte var de kommer ifrån, men de säkert kommer,Jag hoppas att de comin 'för mig!Och jag vet inte hur de gör det, men de säkert göra det bra,Jag hoppas att de doin det gratis!De ger mig cat scratch fever ... cat scratch fever!Första gången som jag fick det jag var bara tio år gammal,Fick det från kitty intill ...Jag gick till doktorn och han gav mig ett botemedel,Jag tror jag fick det lite mer!Fick en dålig repa feber ...
		-- Ted Nugent, "Cat Scratch Fever"

%
Jo, min pappa flyttade hemifrån när jag var tre,Och han inte lämnar mycket för Ma och mig,Bara och gamla gitarr an'a tom flaska sprit.Nu Jag klandrar inte honom för att han sprang och gömde,Men den ringaste sak som han någonsin gjorde,Var innan han lämnade han gick och namngav mig Sue....Men jag gjorde mig ett löfte till månen och stjärnorna,Jag skulle söka honkey tonks och barer,Och döda mannen som ger mig denna fruktansvärda namn.Det var Burg i mitten av juli,Jag skulle bara drabba staden och min hals var torr,Trodde jag skulle sluta och har själv en brygga,Vid en gammal saloon på en gata i lera,Sitter vid ett bord, som handlar stud,Satt det smutsiga (bleep) som namngav mig Sue....Nu visste jag att ormen var min egen söta pappa,Från en wornout bild som min mor hade,Och jag visste att ärr på kinden och hans onda ögat ...
		-- Johnny Cash, "A Boy Named Sue"

%
Jo, min terminalens inlåst, och jag har inte fått någon post,Och jag kan inte minnas den senaste gången mitt program inte misslyckas;Jag har högar i mina structs, jag har arrayer i mina köer,Jag har fått: Segmente brott - Kärn dumpade blues.Om du tycker att det är trevligt att du får vad du C,Gå sedan: ologisk uttalande med hela din familj,"Orsak Högsta domstolen är inte det enda stället med: utsikt bussfel.Jag har fått: Segmente brott - Kärn dumpade blues.På en PDP-11, ska livet vara en vind,Men med VAXen i huset även magnetband skulle frysa.Nu kanske du tror att till skillnad från VAXen jag skulle veta vem jag missbrukar,Jag har fått: Segmente brott - Kärn dumpade blues.
		-- Core Dumped Blues

%
Tja, vissa tar glädje i vagnarna en rullande,Och vissa tar glädje i hurling och bowling,Men jag tar glädje i saften av korn,Och uppvakta ganska rättvist pigor på morgonen ljusa och tidigt.
		-- Core Dumped Blues

%
Tja, vi stora rocksångare, vi har fått gyllene fingrar,Och vi älskade överallt vi gå.Vi sjunger om skönhet, och vi sjunger om sanningen,Vid tio tusen dollar per show.Vi tar alla typer av piller för att ge oss alla typer av spänning,Men spänningen vi har aldrig känt,Är spänningen som kommer get'cha, när du får din bild,På omslaget av Rolling Stone.Jag fick en freaky gammal dam, namn Cole kung Katie,Som broderar på mina jeans.Jag fick min stackars gamla gråhåriga pappa,Drivin min limousine.Nu är det alla utformade för att blåsa våra sinnen,Men våra sinnen kommer inte att verkligen blåsas;Liksom slag som kommer get'cha, när du får din bild,På omslaget av Rolling Stone.Vi fick en massa små, teen-aged, blåögda groupies,Vem gör vad som helst vi säger.Vi fick en äkta indisk guru, som är Inlärning "oss ett bättre sätt.Vi fick alla vänner som pengar kan köpa,Så vi aldrig behöver vara ensam.Och vi fortsätter gettin 'rikare, men vi kan inte få vår bild,På omslaget av Rolling Stone.[Som en anteckning, så småningom de gjorde omslaget till RS. Ed.]
		-- Dr. Hook and the Medicine Show

%
Vad hemskt ironi är detta?Vi är som gudar, men vet att det inte.
		-- Dr. Hook and the Medicine Show

%
Vad gjorde ya göra med din börda och ditt kors?Har du bär den själv eller har du gråta?Du och jag vet att en börda och ett kors,Kan endast utföras på en mans rygg.
		-- Louden Wainwright III

%
Vad händer med en dröm uppskjuten?Är det torka uppSom ett russin i solen?Eller gro som en öm -Och sedan köra?Är det stinker som ruttet kött?Eller skorpa och socker över -Som en sirapsliknande söt?Kanske är det bara bottnarSom en tung last.Eller betyder explodera?
		-- Langston Hughes

%
Vad har rötter som ingen ser,Är högre än träden,Upp, upp det går,Och ändå aldrig växer?
		-- Langston Hughes

%
Vilka smärtor andra njutning mig,Hemma är jag i Lisp eller C;Det i soffan i extas,'Til debugger s peta i fly,I kärnminnet.I systemet utrymme, systemutrymme, ska det i fare--Insidan av en VAX på en kisel kvadrat.
		-- Langston Hughes

%
Vad segmentets detta, att, som att vilaPå FHA0, sover?Vad systemfil, låg här ett tag här, detta är "acct.run"Medan hackare runt det var gråt? Redovisning fil för alla.Dumpa, dumpa det och skriver ut det,Filen är highseg av inloggning.Varför ligger det här, om offentlig diskOch varför är det nu oskyddade?Ett fel i Incant, gjorde det så. Mount, montera alla dina DECtapes nuOch kopiera filen på något sätt, på något sätt. Problemet har inte korrigerats.Dumpa, dumpa det och skriver ut det,Filen är highseg av inloggning.
		-- to Greensleeves

%
Vad vi är Guds gåva till oss.Vad vi Bli är vår gåva till Gud.
		-- to Greensleeves

%
Vad med ChromoDynamics och elektro alltförVår standardiserad modell bör tillfredsställa även dig,Tho "när du sa att charm fanns ingenDet krävdes mod för att växla så att säga jorden rör sig inte Sun.Ändå din State of the Union näst sista storaÄr den sista kända tillhåll för Fractional Charge,Och när du surfar i bubbelpoolen med surdeg rulleVänligen fundera tidens din enda Monopole.Dina OS var roligt, du bör föra dem alla tillbakaFör transsexuell tennis eller Anamalon Track,Men Hollywood-filmer förblir sinfully råaVare sett på teve eller Fjärr Sett.Nu spänn fast sunbelts, för du har gjort det en gång,Du sa det i Leipzig av det vi tillber,Att du har byggt en otrolig kristallin sfärVars tyska skötare spridda darrande och rädslaAv döden av vår teori genom partikel ZetaSom jag ska satsa är inte det säga din artikel, senare.
		-- Sheldon Glashow, Physics Today, December, 1984

%
Vad är kärlek men en andrahands känslor?
		-- Tina Turner

%
Vad lever fortfarande på tjugotvå,En ren upprättstående chap som du?Visst, om din hals "tis svårt att skära,Slits din flicka, och gunga för det.Liksom nog kommer du inte vara glad,När de kommer att hänga dig, lad:Men bacon är inte det endaDet är botas genom att hänga från en sträng.Så när utspillt bläck i nattenSprider o'er blotting dyna av ljus,Lads vars uppgift är fortfarande att göraSka vässa sina knivar, och tänker på dig.
		-- Hugh Kingsmill

%
När ett lejon möter en annan med en högre vrål,den första lion tror den sista en borrning.
		-- G. B. Shaw

%
När jag tänker på mig själv,Jag nästan skrattar ihjäl mig,Mitt liv har varit ett mycket stort skämt, Sextio år i dessa folks världEn dans som är gick Barnet jag fungerar för samtal mig flickaEn låt som är eker, jag säger "Ja frun" för att arbeta skull.Jag skrattar så hårt jag nästan kväva för stolt för att böjaNär jag tänker på mig själv. Alltför dålig för att bryta,Jag skrattar tills min magen,När jag tänker på mig själv.Mina föräldrar kan få mig att dela min sida,Jag skrattade så hårt jag nästan dog,De berättelser de berättar, låter precis som att ligga,De växer frukten,Men äter skalet,Jag skrattar tills jag börjar gråta,När jag tänker på mina föräldrar.
		-- Maya Angelou

%
När i panik, rädsla och tvivel,Dricka i fat, äta, och skrika.
		-- Maya Angelou

%
När i denna värld rubriker läsaAv dem vars hjärtan är fyllda med girighetVem råna och stjäla från dem som behöverRopet går upp med bländande hastighet för Underdog (UNDERLÄGE!)Underdog (UNDERLÄGE!)Blixtens hastighet, bruset av åskaKampen mot alla som råna eller plundringUnderdog (ah-ah-ah-ah)underlägeUNDERLÄGE!
		-- Maya Angelou

%
När de har problem eller tvivel,köra i cirklar, skrika och ropa.
		-- Maya Angelou

%
När licensavgifter är för höga,användare gör saker för hand.När ledningen är alltför påträngande,användare förlorar sin själ.Hack för användarens nytta.Lita på dem; lämna dem ifred.
		-- Maya Angelou

%
När kärleken är borta, det finns alltid rättvisa.Och när rättvisa är borta, det finns alltid kraft.När kraft är borta, det finns alltid mamma.Hej mamma!
		-- Laurie Anderson

%
När mina näve knyter knäcka det öppna,Innan jag använder den och förlorar min cool.När jag ler berätta några dåliga nyheter,Innan jag skrattar och agera som en idiot.Och om jag sväljer något ont,Sätt dig finger ner min hals.Och om jag ryser ge mig en filt,Hålla mig varm låt mig bära din jackaIngen vet hur det är att vara dålig människa,att vara ledsen man.Bakom blåa ögon.Ingen vet hur det är att vara hatad,som skall fated,Att berätta bara ligger.
		-- The Who

%
Då syre Tech spelade Väte U.Spelet hade just börjat när Väte gjorde två snabba poängOch Oxygen hade fortfarande ingenDå Oxygen gjorde ett enda målOch så förblev, vid Väte 2 och syre ettKallad på grund av regn.
		-- The Who

%
När någon gör ett drag Vi skickar dem allt vi har,Som vi inte godkänner, John Wayne och Randolph Scott,Vem är det som alltid ingriper? Kom ihåg de spännande kampscener?FÖRENTA NATIONERNA och O.A.S., till stranden i Tripoli,De har sin plats, antar jag, men inte Mississippoli,Men först, skicka flottorna! Vad gör vi? Vi skickar flottorna!För den starkes rätt, medlemmar av kårenOch tills de har sett ljuset, alla hatar tanken på krig:De måste skyddas, skulle de hellre döda dem genomfredliga medel.Alla sina rättigheter respekterade, Sluta kalla det aggression--Till någon vi vill kan väljas. Vi hatar det uttrycket!Vi vill bara att världen ska vetaAtt vi stöder status quo;De älskar oss överallt vi går,Så när du är osäker, skicka flottorna!
		-- Tom Lehrer, "Send The Marines"

%
När Guru administrerar, användarnaär knappast medveten om att han existerar.Nästa bästa är en sysop som är älskad.Därefter en som fruktas.Och värst, en som föraktas.Om du inte litar på användarna,du gör dem opålitliga.Guru inte prata, han hackar.När hans arbete är gjort,användarna säger, "Amazing:vi genomfört det, alla av oss! "
		-- Tom Lehrer, "Send The Marines"

%
När ledarna talar om fredVanligt folk vetDet kriget kommerNär ledarna förbannar krigetMobiliseringen ordern redan skrivit ut.Varje dag, för att tjäna mitt dagliga brödJag går till marknaden där ligger köpsFörhoppningsvisJag tar min plats bland säljarna.
		-- Bertolt Brecht, "Hollywood"

%
När användarna ser ett GUI så vacker,andra användargränssnitt blir ful.När användarna se vissa program som vinnare,andra program blir lossage.Pekare och NULL referera varandra.Hög nivå och assembler beroende av varandra.Dubbel och flyta gjutna till varandra.Hög endian och låg endian definiera varandra.Tag och tills följa varandra.Därför Guruprogram utan att göra någontingoch undervisar utan att säga något.Varningar uppstår och han låter dem komma;processer byts och han låter dem gå.Han har men inte besitter,fungerar men inte förväntar sig.När hans arbete utförs, raderar han det.Det är därför det varar för evigt.
		-- Bertolt Brecht, "Hollywood"

%
När du och jag är långt ifrån varandraKan sorg bryta ert anbud hjärta?Jag älskar dig älskling, ja jag gör;Sömn är så söt när jag drömmer om dig;Allt du är en blommande ros.Night är här så jag måste stänga.Med omsorg läsa det första ordet av varje rad.Du hittar en fråga till mig.
		-- Yours hopefully, The VAX.

%
När du befinner dig i fara,När du hotas av en främling,När det ser ut som du kommer att ta en lickin '...Det finns en sak du bör lära,När det inte finns någon annan att vända sig till,Caaaall för Super kyckling !! (** Bwuck-bwuck-bwuck-bwuck **)Caaaall för Super kyckling !!
		-- Yours hopefully, The VAX.

%
När du får vad du vill ha i din kamp för självOch världen gör dig till kung för en dag,Bara att gå till en spegel och titta på dig självOch se vad den mannen har att säga.För det är inte din pappa eller mamma eller fruVars dom över dig måste passera;Stipendiaten vars dom räknas mest i ditt livÄr en stirrar tillbaka från glaset.Vissa människor kanske tror att du en rak shootin "kamratOch ringa dig en underbar kille,Men mannen i glaset säger att du är bara en luffareOm du inte kan se honom rakt i ögonen.Han är karl att behaga, strunt alla de andra,För han är med dig klar fram till slutet,Och du har klarat din farligaste, svårt testOm mannen i glaset är din vän.Du kan lura hela världen ner vägen i livetOch få klapp på ryggen när du passerar,Men den slutliga belöningen blir sorger och tårarOm du har lurat mannen i glaset.
		-- Yours hopefully, The VAX.

%
När du möter en mästare krigare,visa honom ditt svärd.När du möter en man som inte är en poet,inte visar honom din dikt.
		-- Rinzai, ninth century Zen master

%
När du overesteem stora hackare,fler användare blir cretins.När du utvecklar kryptering,fler användare blir kex.The Guru ledergenom att tömma användarens sinnenoch öka sina kvoter,genom att försvaga deras ambitionoch hårdare deras beslutsamhet.När användare saknar kunskap och lust,förvaltning kommer inte att försöka ingripa.Öva inte-looping,och allt faller på plats.
		-- Rinzai, ninth century Zen master

%
När du är en JappDu är en Japp hela vägenFrån din första skiva BrieTill din sista Cabernet.När du är en JappDu är inte bara en drömmareDu gör saker att händaDu kör en Beamer.
		-- Rinzai, ninth century Zen master

%
När du är borta, jag är rastlös, ensam,Eländiga, tråkigt, nedslagen; endastHär är där skon klämmer, min älskling kärtJag känner samma när du är nära.
		-- Samuel Hoffenstein, "When You're Away"

%
När Richard Cory gick centrum,Vi människor på trottoaren såg på honom:Han var en gentleman från sula till kronan,Ren gynnade och imperiet smal.Och han var alltid tyst klädd,Och han var alltid mänsklig när han talade;Men han fladdrade pulser när han sade:"God morgon", och han glittrade när han gick.Och han var rik - ja, rikare än en kung -Och beundransvärt skolad i varje nåd:Vid fint, trodde vi att han var alltFör att göra oss önskar att vi var i hans ställe.Så om vi arbetade, och väntade på ljus,Och gick utan kött, och förbannade brödet;Och Richard Cory, en lugn sommarnatt,Gick hem och sätta en kula genom huvudet.
		-- E. A. Robinson, "Richard Cory"

%
VAR KAN ärendetÅh, kära, där kan ärendet varaNär det omvandlas till energi?Det finns en liten förlust av paritet.Johnnys så länge på mässan.
		-- E. A. Robinson, "Richard Cory"

%
Var är mannen kan underlätta ett hjärtaSom en satängkappa?
		-- Dorothy Parker, "The Satin Dress"

%
Där, oh, där är du i kväll?Varför lämnade du mig här ensam?Jag sökte över hela världen, och jag trodde att jag hade hittat den sanna kärleken.Du träffade en annan, och * PPHHHLLLBBBBTTT *, wuz du borta.Gloom, förtvivlan och vånda på mig.Djup mörk depression, överdriven elände.Om det inte vore för otur, skulle jag har ingen tur alls.Åh, dysterhet, förtvivlan och vånda på mig.
		-- Hee Haw

%
Vare sig trötta eller unweary, o människa, inte vila,Upphör inte din ensam kamp.Gå på, inte vila.
		-- An old Gujarati hymn

%
Om du kan höra det eller inte,Universum skrattar bakom ryggen.
		-- National Lampoon, "Deteriorata"

%
Medan Europas öga fix'd på mäktiga saker,Ödet för imperier och hösten kungar;Medan kvacksalvare statliga måste varje producera sin plan,Och även barn läspa rättigheter Man;Mitt i denna mäktiga väsen låt mig nämna,Rätterna av kvinnan förtjänar viss uppmärksamhet.
		-- Robert Burns, Address on "The Rights of Woman", 26/10 1792

%
Medan jag nickade nästan tupplur, plötsligt kom en avlyssning,Som av någon försiktigt rappa, rappa på min kammardörr.[Citerat i "VMS interna och datastrukturer", V4.4, närhänvisning till hårdvaruavbrott.]Och nu ser jag med ögat lugnDen mycket puls av maskinen.[Citerat i "VMS interna och datastrukturer", V4.4, närmed hänvisning till mjukvaru avbrott.]
		-- William Wordsworth, "She Was a Phantom of Delight"

%
Medan promenader ner en fullsattStadsgata häromdagen,Jag hörde en liten sjöborreTill en kamrat vända och säga,"Säg, Chimmey, lemme berätta youse,Jag skulle vara glad som en musslaOm jag bara var de fällare datMig Mudder t'inks jag."Hon t'inks jag ett konstigt, mina vänner, bli din ett liv i slitEn "hon vet sin lilla pojke eller outspädd glädje,Kunde aldrig blanda wit "nuttin" Du kan lära en hälsosam läxaDat var ful, medelvärdet eller dåligt. Från den lilla, untutored pojke.Åh, mycket o gånger jag sitta och t'ink inte sträva efter att vara en jordisk helgonHur trevligt "twould vara, gee vina! Med blicken fäst på en stjärna:Om en fällare var de fällare Försök att vara karl somDat hans mudder t'inks han är. "Din mamma tycker du är.
		-- Will S. Adkin, "If I Only Was the Fellow"

%
Piska, baby.Vispa det rätt.Piska, baby.Vispa det hela natten!
		-- Will S. Adkin, "If I Only Was the Fellow"

%
Vem älskar inte vin, kvinnor och sång,Förblir en dåre hela sitt liv länge.
		-- Johann Heinrich Voss

%
Vem älskar inte klokt men alltför välSer ut på Helen ansikte i helvetet,Men han vars kärlek är tunn och visKommer att betrakta John Knox i paradiset.
		-- Dorothy Parker

%
Vem gjorde världen jag kan inte säga;'Tis gjort, och här är jag i helvetet.Min hand, men nu knogarna blöder,Jag har aldrig nedsmutsade med en sådan handling.
		-- A. E. Housman

%
Vem ska själv är lag inget lag doth behovkränker ingen lag, och är en kung faktiskt.
		-- George Chapman

%
Varför tittar du påTvättmaskinen?Jag älskar underhållningSå länge det är ren.Professor Doberman:Medan föregående dikt är onekligen en förändring från bevakadepessimism "The Hound of Heaven," det kan inte betraktas som en okvalificeradförbättring. Grumlighet är av värde endast då det tenderar att klargöra poetiskaerfarenhet. Så mycket som en tvingas att beundra diktens teknik, enmåste ifrågasätta huruvida dess byplay av komplexa litterära allusioner inte iFaktum distrahera från enheten i det hela. I den slutliga analysen, enfår en stark känsla av att dikten längd kunde säkert hareducerats med en faktor av åtta eller tio utan att offra något av dessmenande. Det är önskvärt att ytterligare offentliggörandet av denna dikt kan varaavvaktan en grundlig undersökning av dess potentiella subversivakonsekvenser.
		-- George Chapman

%
Med / Utan - och som kommer att förneka det är vad striderna all om?
		-- Pink Floyd

%
Vaknade upp denna mornin 'en' Jag hade själv en öl,Ja, Ah vaknade i morse "en" Jag hade själv en ölFramtiden osäkra och slutet är alltid nära.
		-- Jim Morrison, "Roadhouse Blues"

%
Vaknade i morse, inte tro vad jag såg.Hundra miljarder flaskor spolas upp på stranden.Verkar jag inte ensam om att vara ensam.Hundra miljarder skeppsbrutna söker ett samtal.
		-- The Police, "Message in a Bottle"

%
Ja från bordet av mitt minneJag ska torka bort alla triviala förtjust poster.
		-- Hamlet

%
Ja mig, jag fick en flaska framför mig.Och Jimmy har en frontal lobotomi.Bara olika sätt att döda smärtan densamma.Men jag vill hellre ha en flaska framför mig,Än att ha att ha en frontal lobotomi.Jag kan drickas men åtminstone jag inte galen.
		-- Randy Ansley M.D. (Dr. Rock)

%
Igår på den trappJag träffade en man som inte var där.Han var inte där i dag igen -Jag tror att han är från CIA.
		-- Randy Ansley M.D. (Dr. Rock)

%
"Du är gammal, fadern William" den unge mannen sade,"Alla dina papper dessa dagar ser likadana;De Williams skulle vara bättre oläst -Har dessa fakta fylla dig aldrig med skam? ""I min ungdom," Fader William svarade till sin son,"Jag skrev underbart papper i överflöd;Men den stora rykte jag upptäckte att jag hade vunnit,Gjorde det meningslöst att tänka längre. "
		-- Randy Ansley M.D. (Dr. Rock)

%
"Du är gammal, far William," den unge mannen sade,"Och håret har blivit mycket vitt;Och ändå ständigt stå på huvudet -Tror du på din ålder, är det rätt? ""I min ungdom", svarade pappa William till sin son,"Jag fruktade det kan skada hjärnan;Men nu när jag är helt säker har jag ingen,Varför gör jag det igen och igen. ""Du är gammal", sa ynglingen ", som jag nämnde tidigare,Och har vuxit mest ovanligt fett;Men du vände en back-kullerbytta in genom dörren -Be vad är orsaken till det? ""I min ungdom," sade den vise, när han skakade grå lås,"Jag höll alla mina lemmar mycket smidigGenom användning av denna salva - en shilling lådan -Tillåt mig att sälja dig ett par? "
		-- Randy Ansley M.D. (Dr. Rock)

%
"Du är gammal", sade ungdom "och jag har fått veta av mina kamraterAtt dina föreläsningar bar människor till döden.Men du prata hundra konventioner per år -Tror du inte att du ska spara din andedräkt? ""Jag har svarat tre frågor och som är tillräckligt"Sade fadern, "Ge inte dig själv luftar!Tror du att jag kan lyssna hela dagen för att sådana saker?Var bort, eller jag ska sparka dig nere! "
		-- Randy Ansley M.D. (Dr. Rock)

%
"Du är gammal", sade ungdom "och käkarna är för svagFör något hårdare än talg;Men du avslutade gås, med ben och näbb -Be, hur lyckades du göra det? ""I min ungdom," sade fadern, "Jag tog till lagen,Och hävdade varje fall med min fru;Och muskelstyrka som det gav till min käke,Har varat resten av mitt liv. ""Du är gammal", sade ungdom "skulle knappast troAtt ögat var så stabil som någonsin;Men du balanserad en ål på slutet av näsan -Vad gjorde du så väldigt smart? ""Jag har svarat tre frågor, och det är tillräckligt"Sade fadern. "Ge inte dig själv airs!Tror du att jag kan lyssna hela dagen för att sådana saker?Var bort, eller jag ska sparka dig nedför trappor! "
		-- Randy Ansley M.D. (Dr. Rock)

%
"Du är gammal", sade ungdom "och dina program körs inte,Och det finns inte ett språk du vill,Ändå av användbara förslag om hjälp du har ingen -Har du funderat på att ta en vandring? ""Eftersom jag aldrig skriva program", hans far svarade,"Varje språk ser lika illa;Ändå människor fortsätta att betala för att läsa alla mina böckerOch inser inte att de har haft. "
		-- Randy Ansley M.D. (Dr. Rock)

%
"Du är gammal", sa ynglingen ", som jag nämnde tidigare,Och göra fel fåtal personer kan bära;Du klagar allas engelska men er -Tror du verkligen att detta är ganska rättvist? ""Jag gör massor av misstag," Fader William förklarade,"Men min resning i dessa dagar är så storAtt ingen kritiker kan skada mig - Jag har dem alla rädda,Och för att stoppa mig är det nu alldeles för sent. "
		-- Randy Ansley M.D. (Dr. Rock)

%
Du kan kräla med en älskare, du kan kräla med en vän,Du kan kräla med din chef, och det har aldrig ta slut.(Kör) Grovel, kräla, kräla, varje natt och varje dag,Kräla, krypa, kräla i din egen märkliga sätt.Du kan krypa i en hall, kan du kräla i en park,Du kan krypa i en gränd med en rånare after dark.(kör)Du kan kräla med din farbror, du kan kräla med din faster,Du kan kräla med Apple, även om du säger att du inte kan.(kör)
		-- Randy Ansley M.D. (Dr. Rock)

%
Du går ner till pickup stationen,sugen värme och skönhet;Du nöja sig med mindre än fascination -några drinkar senare du inte är så kräsen.Och de sista lamporna strippa skuggornapå denna märkliga nya kött du har hittat -Kramade natten till dig som ett fikonlövdu skynda till svärtanoch filtar att fastställa ett intryckoch din ensamhet.
		-- Joni Mitchell

%
Du måste betala dina skulder om du vill sjunga blues,Och du vet att det inte kommer lätt ...Jag inte begära för mycket, jag vill bara förtroende,Och du vet att det inte kommer lätt ...
		-- Joni Mitchell

%
Du vet mitt hjärta håller tellin "mig,Du är inte en unge på trettiotre,Du spelar runt du förlorar din fru,Du spelar för länge, förlorar du ditt liv.Några mĺste vinna, några mĺste förlora,Goodtime Charlies fick blues.
		-- Joni Mitchell

%
Du kan vara rätt, jag kan vara galen,Men det bara kan vara en galning du letar efter!
		-- Billy Joel

%
Du hittar mig dricka ginI den lägsta typ av inn,Eftersom jag är en stel Vegetariskt.
		-- G. K. Chesterton

%
Du kommer alltid att vara,Vad du alltid var,Som inte har någonting att göra med,Allt för att göra, med henne.
		-- Company

%
Dina vise män vet inte hur det kännsAtt vara tjock som en tegelsten.
		-- Jethro Tull, "Thick As A Brick"

%
Ers Nåd är dina ugnarsom i likhet med gamla idoler, förlorade obscenes,har smält tarmarna; din vision ärmaskiner för tillverkning av flera maskiner.
		-- Gordon Bottomley, 1874

%
Yours är inte anledningen,Bara för att Sail Away.Och när du upptäcker att du måste kastaDin Legacy bort;Kom ihåg liv som var det är,Och är så att säga;Chasing ljud över hela galaxen"Till tystnad är bara en oskärpa.
		-- QYX.

%
Vi hittade dig gömmerVi hittade dig liggandeKvävning på smuts och sand.Dina tidigare härligheterOch alla berättelserDras och tvättades med ivriga händer.
		-- ``Cities in Dust'', "Tinderbox", Siouxsie & the Banshees.

%
