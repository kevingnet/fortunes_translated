1893 Den idealiska hjärnan tonic1900 dryck Coca-Cola - läcker och uppfriskande - 5 cent allssoda fontäner1905 Är favoritdryck för damer när törstiga - trött - förtvivlad1905 Uppdaterar trötta, ljusare intellekt och rensar hjärnan1906 Drycken kvalitets1907 Bra till sista droppen1907 Den uppfyller törst och behagar gommen1907 uppfriskande som en sommarbris. Förtjusande som ett dopp i havet1908 dryck som Cheers men inte BERUSA1917 Det finns en läcker friskhet i smaken av Coca-Cola1919 Det uppfyller törst1919 Smaken är testet1922 Varje glas har svaret på törst1922 Törst vet ingen säsong1925 Njut av sällskaplig drink
		-- Coca-Cola slogans

%
1925 med en drink så bra, 'tis dårskap att vara törstig1929 Den höga tecken på förfriskningar1929 Pausen som uppdateras1930 Det skulle vara bra att få där det är1932 Drycken som gör en paus uppfriskande1935 Pausen som ger vänner tillsammans1937 stopp för en paus ... GO uppdateras1938 Den bästa vän törst någonsin haft1939 Törst slutar här1942 Det är the real thing1947 Ha en cola1961 Zing! Vilken uppfriskande ny känsla1963 Saker går bättre med koks1969 Face Uncle Sam med en cola i handen1979 Ha en cola och ett leende1982 Koks är det!
		-- Coca-Cola slogans

%
Ett par av barnen försökt med pickles i stället för paddlar för en Ping-Pongspel. De hade volley av Dills.
		-- Coca-Cola slogans

%
En gård på landet hade flera kalkoner, var det känt somhus av sju slukar.
		-- Coca-Cola slogans

%
En gourmet som tänker på kalorier är som en tårta som ser på klockan.
		-- James Beard

%
En ny kock från Indien fick sparken en vecka efter att ha startat jobbet. hanhålls gynna curry.
		-- James Beard

%
En midja är en fruktansvärd sak att tänka på.
		-- Ziggy

%
En fru började betjäna hackat kött, måndag hamburgare, tisdag köttlimpa, onsdag tartar biff och torsdag köttbullar. På fredag ​​morgon henneman morrade, "Hur nu, mark ko?"
		-- Ziggy

%
Skådespelare: Så vad gör du för en levande?Doris: Jag arbetar för ett företag som gör bedrägligt grunt serveringrätter för kinesiska restauranger.
		-- Woody Allen, "Without Feathers"

%
Egentligen är mitt mål att ha en smörgås uppkallad efter mig.
		-- Woody Allen, "Without Feathers"

%
"Och vad ska du göra när du växa upp och bli lika stor som mig?"frågade far till sin lilla son."Diet".
		-- Woody Allen, "Without Feathers"

%
Allt är bra om den är gjord av choklad.
		-- Woody Allen, "Without Feathers"

%
Allt som är bra och användbar är gjord av choklad.
		-- Woody Allen, "Without Feathers"

%
När han hade fruktat, hade hans order glömts bort och alla hade förtpotatissallad.
		-- Woody Allen, "Without Feathers"

%
Som med de flesta fina saker, har choklad sin säsong. Det finns en enkelminneshjälp som du kan använda för att avgöra om det är rätt tidatt beställa choklad rätter: varje månad vars namn innehåller bokstaven A,E, eller U är den rätta tidpunkten för choklad.
		-- Sandra Boynton, "Chocolate: The Consuming Passion"

%
Var försiktig när du bita i din hamburgare.
		-- Derek Bok

%
BUA! Vi ändrade Coke igen! BLEAH! BLEAH!
		-- Derek Bok

%
Bojkott kött - suga tummen.
		-- Derek Bok

%
Carob fungerar enligt principen att när de blandas med rätt kombination avfett och socker, kan det duplicera choklad i färg och konsistens. Självklart,samma kan sägas om smuts.
		-- Derek Bok

%
Ost - mjölk språng mot odödlighet.
		-- Clifton Fadiman, "Any Number Can Play"

%
Kinesiskt talesätt: "Han som talar med kluven tunga, inte behöver ätpinnar."
		-- Clifton Fadiman, "Any Number Can Play"

%
Tänk på följande axiom noga:"Allt är bättre när det sitter på en Ritz."och"Allt är bättre med Blue Bonnet på det."Vad händer om man sprider Blue Bonnet margarin på en Ritz smällare? DeTanken är skrämmande. Är detta hur Gud kom till? Försök att inteöverväga det faktum att "Saker går bättre med koks".
		-- Clifton Fadiman, "Any Number Can Play"

%
Kära Mister Språk Person: Jag är nyfiken på uttrycket, "En del avDetta komplett frukost ". Hur det kommer upp är, min 5-åriga varatittar på TV tecknad visar på morgonen, och de kommer att visa en reklamfilm förbarn komprimerad frukost förening såsom "Froot Loops" eller "TurCharms ", och de visar alltid det sitter på ett bord bredvid några faktiska matsåsom ägg, och speakern alltid säger: "En del av denna fullständigaFrukost ". Inte som verkligen betyder," I anslutning till detta komplett frukost ",eller "På samma bord som denna komplett frukost"? Och kunde de inte göraväsentligen samma krav om man istället för Froot slingor, sätter de en burkrakkräm där, eller en död fladdermus?Svar: Ja.
		-- Dave Barry, "Tips for Writer's"

%
Död före vanära. Men varken före frukost.
		-- Dave Barry, "Tips for Writer's"

%
Hörde du att kapten Crunch, Sugar Bear, Tony Tiger, ochSnap, Crackle och Pop var alla mördades nyligen ...Polisen misstänker att arbetet i en spannmåls mördare!
		-- Dave Barry, "Tips for Writer's"

%
Dieters leva livet i fasta lane.
		-- Dave Barry, "Tips for Writer's"

%
Middagen är klar när röken larmet utlöses.
		-- Dave Barry, "Tips for Writer's"

%
Dricker inte kaffe i början av A.M. Det kommer att hålla dig vaken fram till middagstid.
		-- Dave Barry, "Tips for Writer's"

%
Oroa dig inte om vilken sida brödet är smörade på: du äter båda sidor.
		-- Dave Barry, "Tips for Writer's"

%
Känner du personligen ansvarig för världslivsmedelsbristen?Varje gång du går till stranden, inte på strömmen komma in?Har du någonsin ätit en hel älg?Kan du se din hals?Gör joggare ta varv runt dig för motion?Om så är fallet, välkommen till National Fat vecka.Den här veckan ska vi äta utan skuld, och kick off vår kampanj för medlemskap,... Genom tvångsmatning en låda av majsstärkelse till en mager person.
		-- Garfield

%
Under den amerikanska revolutionen, en britt försökte plundra en gård. hansnubblat över en sten på marken och föll, varpå en aggressiv RhodeIsland Red hoppade på toppen. Att se detta bonden kommenterade, "Chicken catchen Tory! "
		-- Garfield

%
Ät så mycket du vill - bara inte svälja det.
		-- Harry Secombe's diet

%
Äta dricka och vara glada! Tommorrow du kan vara i Utah.
		-- Harry Secombe's diet

%
Äta dricka och vara glada, för i morgon kan de göra det olagligt.
		-- Harry Secombe's diet

%
Äta dricka och vara glada, ty i morgon vi diet.
		-- Harry Secombe's diet

%
Äta rätt, hålla formen, och dö i alla fall.
		-- Harry Secombe's diet

%
"Ät, drick och var glad, för i morgon kan du arbeta."
		-- Harry Secombe's diet

%
Äta choklad är som att vara kär utan försämringen.
		-- Harry Secombe's diet

%
Även en blind gris snubblar på några ekollon.
		-- Harry Secombe's diet

%
Även en kål kan titta på en kung.
		-- Harry Secombe's diet

%
Varje gång jag gå ner i vikt, finner det mig igen!
		-- Harry Secombe's diet

%
Allt jag är antingen olagligt, omoraliskt eller gödning.
		-- Alexander Woollcott

%
Allt är värt exakt lika mycket som en rapa, varvid skillnaden äratt en rapa är mer tillfredsställande.
		-- Ingmar Bergman

%
Fett Liberation: eftersom en midja är en fruktansvärd sak att tänka på.
		-- Ingmar Bergman

%
Feta människor i världen förenar, har vi inget att förlora!
		-- Ingmar Bergman

%
Tankeställare är inget substitut för the real thing.
		-- Walt Kelly, "Potluck Pogo"

%
För er som har varit olyckligt nog att aldrig har smakat"Stor Chieftain O 'Pudden Race" (dvs haggis) här är ett lätt att följarecept som resulterar i en maträtt anmärkningsvärt lik den ovan nämndaskyddade arter.ingredienser:En fåra Pluck (hjärta, lungor, lever) och väska2 teacupsful rostade havregryn1 tesked salt8 oz. strimlad talg2 små lökar1/2 tesked svartpepparSkrapa och ren väska i kallt, sedan varmt vatten. Blötlägg i saltvattenöver natten. Tvätta mod, sedan koka i 2 timmar med luftstrupen dränering överden sida av potten. Behålla en pint lager. Skär av luftstrupen, ta bort överskottbrosk, hacka eller färs hjärta och lungor, och riv bästa delen av levern (omendast hälften). Förvälla och hacka lök, blanda tillsammans med havregryn, talg,salt, peppar och lager för att fukta. Packa blandningen i påsen, vilket möjliggörsvullnad. Koka i tre timmar, stickande regelbundet överallt. Om påsen intetillgängliga, ånga i smord bassäng omfattas av smörpapper och tyg förfyra till fem timmar.
		-- Walt Kelly, "Potluck Pogo"

%
Fortune Bidrag från månad till Djurrätts Debatt:Jag ska hålla sig borta från djurens sätt om de ska hålla sig borta från gruvan."Hej du, gå av min tallrik"
		-- Roger Midnight

%
Fortune kost sanningar:1: Glöm vad kokböcker säga, smakar vanlig yoghurt ingenting som gräddfil.2: Alla recept kräver sojabönor smakar lera.3: Carob är inte en godtagbar ersättning för choklad. I själva verket är inte carob    en godtagbar ersättning för något, utom kanske brun skokräm.4: Det finns något sådant som en "kul sallad." Så låt oss sluta låtsas och se    sallader för vad de är: Guds straff för att vara fett.5: Fruktsallad utan maraschino körsbär och marshmallows är ungefär lika    talande som ljummet öl.6: En värld saknar sås är en tragisk plats!7: Du bör omedelbart skicka upp några recept med titeln "läcker och    låg-cal. "Också hoppa rätter med" levande lever. "De är inte och    det inte är.8: Iklädd en ögonbindel ofta gör att många kost livsmedel mer tilltalande.9: Färsk frukt är inte dessert. Kakan är dessert!10: Okra smakar något sämre än namnet antyder.11: En vanlig bakad potatis är inte värt ansträngningen inblandade i tugga och    svälja.
		-- Roger Midnight

%
Gud måste ha älskat kalorier, hon gjorde så många av dem.
		-- Roger Midnight

%
STORA ögonblick i historien (# 7): November 23, 1915Pannkaka smink uppfinns; de flesta människor fortsätter att föredra sirap.
		-- Roger Midnight

%
Har någon någonsin smakade en "slut"? Är de verkligen bitter?
		-- Roger Midnight

%
Har din familj försökt dem?POWDERMILK BISCUITSHeavens, de är välsmakande och snabbt!De är gjorda av fullkornsvete, för att ge blyga personerstyrkan att gå upp och göra vad som behöver göras.POWDERMILK BISCUITSKöpa dem färdiga i den stora blå låda med bilden avkexet på framsidan, eller i den bruna påsen med den mörkafläckar som indikerar friskhet.
		-- Roger Midnight

%
Har en taco.
		-- P. S. Beagle

%
Hem på Range skrevs ursprungligen på nötkött platt.
		-- P. S. Beagle

%
Hors d'oeuvres - en skinksmörgås skuren i fyrtio stycken.
		-- Jack Benny

%
"Hur fick du spendera helgen?" frågade söt brunett sekreterareav sin blonda följeslagare."Fiske genom isen", svarade hon."Fiske genom isen? Vad för?""Oliver."
		-- Jack Benny

%
Hur många hors d'oeuvres är det tillåtet att ta bort en bricka som bärs aven servitör på en trevlig fest?Två, men det finns vägar runt det, beroende på vilken typ av horsd'oeuvre. Om de är de små bakverk saker där du inte kan berätta vad som ärinuti, du tar en, bita av ungefär två tredjedelar av det, sedan säga: "Detta ärost! Jag hatar ost! "Då du lägger resten av det tillbaka på brickan ochbita en annan och gå, "Darn det! En annan ost!" och så vidare.
		-- Dave Barry, "The Stuff of Etiquette"

%
Jag är så optimistisk om priserna på nötkött som jag har just leasade en grytstekmed en option att köpa.
		-- Dave Barry, "The Stuff of Etiquette"

%
Jag bromsar för chezlogs!
		-- Dave Barry, "The Stuff of Etiquette"

%
Jag kunde inte komma ihåg när jag hade varit så besviken. Utom kansketid jag fick reda på att M & Ms verkligen smälter i handen.
		-- Peter Oakley

%
Jag bryr mig inte om socker smakar kommersiella. Jag tycker inte om tanken påen groda hoppar på min frukost.
		-- Lowell, Chicago Reader 10/15/82

%
Jag bryr mig inte där jag sitter så länge jag får utfodras.
		-- Calvin Trillin

%
Jag vet inte ens smör mitt bröd. Jag anser att matlagning.
		-- Katherine Cebrian

%
Jag har inte en ätstörning. Jag äter. Jag får fett. Jag köper nya kläder.Inga problem.
		-- Katherine Cebrian

%
"Jag tycker inte om spenat, och jag är glad att jag inte gör det, för om jag gillade det skulle jagäta det, och jag hatar bara det. "
		-- Clarence Darrow

%
Jag har aldrig varit en att offra min aptit på altaret av utseendet.
		-- A. M. Readyhough

%
Jag har inga tvivel om att det är en del av ödet för den mänskliga rasen,i dess gradvisa förbättringar för att lämna att äta djur.
		-- Thoreau

%
Jag åt bara ett helt paket av söta tårtor och en burk av koks. Jag tror jag såg Gud.
		-- B. Hathrume Duk

%
Jag har aldrig träffat en bit choklad som jag inte gillar.
		-- B. Hathrume Duk

%
Jag aldrig ber före måltid - min mamma är en bra kock.
		-- B. Hathrume Duk

%
"Jag trodde att du försökte komma i form.""Jag är. Formen Jag har valt är en triangel."
		-- B. Hathrume Duk

%
Jag är hungrig, tid att äta lunch.
		-- B. Hathrume Duk

%
Jag har varit på en diet för två veckor och allt jag har förlorat är två veckor.
		-- Totie Fields

%
Om först du fricasee, yngel, stek igen.
		-- Totie Fields

%
Om maten vara musik kärlek, äta upp, äta upp.
		-- Totie Fields

%
Om vitsar var deli kött, skulle detta vara wurst.
		-- Totie Fields

%
Om du är vad du äter, betyder det Euell Gibbons verkligen var en mutter?
		-- Totie Fields

%
Om du placerar din kvällsmat maträtt till örat kan du höra ljudet av enrestaurang.
		-- Snoopy

%
Om du ser en lök ring - besvara den!
		-- Snoopy

%
Om du gryta äpplen som tranbär, de smakar mer som katrinplommon änrabarber gör.
		-- Groucho Marx

%
Om du slösa din tid matlagning, ska du inte missa nästa måltid.
		-- Groucho Marx

%
Om du ska till Amerika, föra din egen mat.
		-- Fran Lebowitz, "Social Studies"

%
Om ditt bröd är inaktuella, göra toast.
		-- Fran Lebowitz, "Social Studies"

%
I Mexiko har vi ett ord för sushi: bete.
		-- Josi Simon

%
Finns det liv innan frukost?
		-- Josi Simon

%
Det är en hård materia, att mina landsmän, argumentera med magen,eftersom den har inga öron.
		-- Marcus Porcius Cato

%
Det gör mig arg när jag går till alla besväret att behöva Marta koka upp omhundra trumpinnar, sedan killen på Marine säger: "Du kan inte kastaatt kyckling till delfinerna. De äter fisk. "Visst de äter fisk om det är allt du ger dem! Man, visa upp.
		-- Jack Handey, The New Mexican, 1988.

%
Det var en modig man som åt den första ostron.
		-- Jack Handey, The New Mexican, 1988.

%
Det skulle vara trevligt om Food and Drug Administration slutade utfärda varningarom giftiga ämnen och bara gav mig namnen på en eller två saker fortfarandesäker att äta.
		-- Robert Fuoss

%
Det är russin som gör inlägg Raisin Bran så raisiny ...
		-- Robert Fuoss

%
Det är så vackert arrangerade på plattan - du vet någons fingrarhar varit över det hela.
		-- Julia Child on nouvelle cuisine.

%
Bara ett fåtal av de perfekta ursäkter för att ha några jordgubbsmousse.Välj en.(1) Det är mindre kalorier än två bitar av jordgubbsmousse.(2) Det är billigare än att gå till Frankrike.(3) Det neutraliserar brownies jag hade igår.(4) Livet är kort.(5) Det är någons födelsedag. Jag vill inte att de fira ensam.(6) Den matchar mina ögon.(7) som sa, "Låt dem äta tårta." måste ha varit att prata med mig.(8) För att straffa mig för att äta dessert igår.(9) Ersättning för all den tid jag tillbringar i duschen inte äta.(10) Strawberry Shortcake är ond. Jag måste hjälpa till att befria världen av det.(11) Jag får svag från att äta allt det friska grejer.(12) Det är den andra årsdagen av natten jag åt vanlig broccoli.
		-- Julia Child on nouvelle cuisine.

%
Killing kalkoner orsakar vintern.
		-- Julia Child on nouvelle cuisine.

%
Kyssa varar inte, matlagning gör.
		-- George Meredith

%
Kök aktivitet är markerad. Smör upp en vän.
		-- George Meredith

%
I natt drömde jag jag åt en tio pund marshmallow, och när jag vaknade uppkudden var borta.
		-- Tommy Cooper

%
Förra veckans husdjur, denna veckas speciell.
		-- Tommy Cooper

%
Låt inte sand i tid få din lunch.
		-- Tommy Cooper

%
Livet är som en skål med soppa med hår flyter på den. Du måsteäta det ändå.
		-- Flaubert

%
"Livet är som en buffé, det är inte bra, men det finns gott om det."
		-- Flaubert

%
Livet är som en burk sardiner. Vi är alla oss, letar efter nyckeln.
		-- Beyond the Fringe

%
Livet är som ett ägg fläck på hakan - du kan slicka det, men det är fortfarandekommer inte att försvinna.
		-- Beyond the Fringe

%
Livet är som en lök: du skal bort det ett lager i taget, och iblanddu gråter.
		-- Carl Sandburg

%
Livet är som en lök: du dra av lager efter lager och sedan hittaDet finns ingenting i det.
		-- James Huneker

%
Livet är för kort för att stoppa en svamp.
		-- Storm Jameson

%
Ett liv utan koffein är stimulerande nog.
		-- Sanka Ad

%
Bor här i Rio, jag har massor av kaffe att välja mellan. Och närdu är på rymmen som jag, uppskattar du en god kopp kaffe.
		-- "Great Train Robber" Ronald Biggs' coffee commercial

%
Hummer:Alla älskar dessa läckra skaldjur, men många kockar ärblödiga om att placera dem i kokande vatten vid liv, som är den endalämplig metod för framställning av dessa. Ärligt talat, det enklaste sättet att eliminera dinskuld är att etablera deras genom att sätta dem på prov innan de tillagas.Faktum är, hummer är bland de mest våldsamma rovdjur på havetgolv, och du bidra till att minska brottsligheten i reven. Ta tag hummerbakom huvudet, ser det rätt i sina otvetydigt skyldiga eyestalks och säga,"Var var du på natten av 21?", Sedan blomstra en bild av enpilgrimsmussla eller en sula och rop, "Kanske kommer detta att uppdatera det råa neuralaapparat du ringer ett minne! "Hummer kommer att våndas märkbart. Det kanäven ta en slägga på dig med en av sina klor. Oförbätterlig. Pop ingrytan. Rättvisa har delgivits, och kort du och dina vänner kommervara också.Husgeråd till ursäkter och ursäkter "
		-- Dave Barry, "Cooking: The Art of Using Appliances and

%
Mannen som anländer till fest två timmar försenat hittar han har blivit slagentill stansen.
		-- Dave Barry, "Cooking: The Art of Using Appliances and

%
MOCK ÄPPELPAJ (behövs ingen äpplen)  Konditorivaror till två crust 9-tums pie 36 Ritz crackers2 dl vatten 2 koppar socker2 tsk grädde av vinsten 2 msk citronsaft  Rivet skal av en citron smör eller margarin  KanelKavla ut botten skorpa bakverk och passar in i 9-tums pajform. Ha sönderRitz crackers grovt i konditorivaror fodrade platta. Kombinera vatten, sockeroch renad vinsten i kastrull, koka försiktigt i 15 minuter. Lägg citronsaft och skal. Häftigt. Häll denna sirap över Crackers, dot generöstmed smör eller margarin och strö kanel. Täck med toppenskorpa. Trim och flöjt kanterna tillsammans. Skär slitsar i topp skorpa att låtaånga fly. Baka i en varm ugn (425 F) 30 till 35 minuter, tills skorpanär skarp och gyllene. Servera varm. Skär i sex till åtta skivor.
		-- Found lurking on a Ritz Crackers box

%
De flesta människor äter som om de gödning sig för marknaden.
		-- E. W. Howe

%
Mountain Dew och munkar ... eftersom frukost är den viktigaste måltidenav dagen.
		-- E. W. Howe

%
Min läkare berättade för mig att sluta ha intima middagar för fyra. Om det inte finnsär tre andra personer.
		-- Orson Welles

%
Min favorit sandwich är jordnötssmör, struntprat, cheddarost, salladoch majonnäs på rostat bröd med ketchup på sidan.
		-- Senator Hubert Humphrey

%
Min vikt är perfekt för min längd - som varierar.
		-- Senator Hubert Humphrey

%
dricker aldrig koks i en rörlig hiss. Hissens rörelse i kombination medkemikalierna i koks producera hallucinationer. Människor tenderar att byta tillödlor och attack utan varning, och stora fladdermöss flyger vanligen ifönster. Dessutom, börjar du tro att hissar har fönster.
		-- Senator Hubert Humphrey

%
äter aldrig något större än ditt huvud.
		-- Senator Hubert Humphrey

%
Aldrig äta mer än du kan lyfta.
		-- Miss Piggy

%
Ingen människa i världen har mer mod än den man som kan stoppa efteräta en jordnöt.
		-- Channing Pollock

%
Ingenting tar smak av jordnötssmör riktigt gillar obesvarad kärlek.
		-- Charlie Brown

%
Nu när du har läst Fortune diet sanningar, kommer du vara beredd på nästagång någon hemmafru eller boutique-ägare som blev kost expert visas på TVatt ansluta sin senaste bok. Och om du fortfarande känner ett styng av skuld föräta kaffe kaka medan du lyssnar på hennes uppmaningar, fråga dig självföljande frågor:(1) Vågar jag lita på en person som faktiskt anser alfalfagroddar enmat?(2) Var författarens enda motiv i att skriva denna bok att bli rikutnyttja övergivna förhoppningar om knubbig människor som mig?(3) Skulle en längre livslängd vara värt om det hade att leva somföreskrivna ... utan fransk friterade lökringar, pizza meddubbel ost, eller enstaka Mai-Tai? (Kom ihåg att levarätt egentligen inte göra dig leva längre, det bara * verkar * somlängre.)Det, och en annan bit av kaffe kaka, borde göra susen.
		-- Charlie Brown

%
jordnöts Blossoms4 koppar socker 16 msk. mjölk4 koppar farinsocker 4 tsk. vanilj4 koppar förkortar 14 koppar mjöl8 ägg 4 tsk. soda4 koppar jordnötssmör 4 tsk. salt-Forma degen till bollar. Rulla i socker och baka på ungreased kakaark vid 375 F. 10-12 minuter. Omedelbart toppen varje kaka med enHersheys kyss eller stjärna trycka ner ordentligt för att knäcka cookie. gör enfan av en hel del.
		-- Charlie Brown

%
Pete: Servitör, är detta kött dåligt.Servitör: Vem har sagt?Pete: Lite svälja.
		-- Charlie Brown

%
Peters hungrig, tid att äta lunch.
		-- Charlie Brown

%
Syltdjurliv - pickle en ekorre idag!
		-- Charlie Brown

%
Katrinplommon ger dig en springa för dina pengar.
		-- Charlie Brown

%
Sätt en kastrull med chili på spisen för att sjuda. Låt det sjuda. Under tiden,halstra en god biff. Äta stek. Låt chili sjuda. Ignorera det.Texas.
		-- Recipe for chili from Allan Shrivers, former governor

%
Sätt katter i kaffet och möss i te!
		-- Recipe for chili from Allan Shrivers, former governor

%
Kom ihåg att DESSERT stavas med två `S medan DESERT stavas meden, eftersom alla vill två desserter, men ingen vill två öknar.
		-- Miss Oglethorp, Gr. 5, PS. 59

%
REGLER FÖR ÄTA - BRONXEN dieter CREED(1) äter aldrig på fastande mage.(2) Lämna aldrig tabellen hungriga.(3) När du reser, aldrig lämna ett land hungrig.(4) Njut av din mat.(5) Njut av din följeslagare mat.(6) verkligen smaka maten. Det kan ta flera portioner tillåstadkomma detta, särskilt om subtilt kryddat.(7) Verkligen känna din mat. Struktur är viktig. Jämföra,till exempel, texturen hos en kålrot med den hos enbrownie. Vilket känns bättre mot dina kinder?(8) äter aldrig mellan snacks, såvida det inte är en måltid.(9) inte känner att du måste avsluta allt på din tallrik. Dukan alltid äta det senare.(10) Undvik vin med ett barnsäkert lock.(11) Undvik blå mat.
		-- Richard Smith, "The Bronx Diet"

%
Heliga kor gör stora hamburgare.
		-- Richard Smith, "The Bronx Diet"

%
Spara gas, inte äta bönor.
		-- Richard Smith, "The Bronx Diet"

%
Ser är lura. Det äter som är tro.
		-- James Thurber

%
Så mycket mat; så lite tid!
		-- James Thurber

%
Vissa indicier är mycket stark, så när du hittar en öring imjölken.
		-- Thoreau

%
Den grundläggande menyalternativ, faktiskt den enda menyalternativet skulle vara ett livsmedel enhet som kallasden "patty", bestående av - skulle garanteras skriftlig - "100procent animaliskt material av något slag. "Alla biffar skulle värmas upp och sedankyls ner i elektroniska apparater omedelbart före servering. DeFrukost Patty skulle vara en bulle på en bulle med sallad, tomat, lök, ägg,Ba-Ko-Bits, Cheez Whiz, en speciell sås gjord genom att hälla ketchup ur enflaska och en liten papperslapp som anger: "Kontrollerad efter nummer 12." DeLunch eller middag Patty skulle vara någon frukost Patties som inte får säljas imorgonen. Seafood Lovers Patty skulle finnas några biffar som varbörjar avge en allvarlig arom. Biffar som också var rank även att varaSkaldjur Lovers Patties skulle pressas till tussar och säljs som "Nuggets."
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Den svarta björnen brukade vara en av de vanligaste sett stora djureftersom i Yosemite och Sequoia nationalparker de bodde utanför av soporoch turistouts. Denna björn har lärt sig att öppna bildörrarna iYosemite, där skador på bilar som orsakas av björnar går till tiotalstusentals dollar om året. Kampanjer för att bearproof alla soporbehållare i vilda områden har varit svårt, eftersom som en biologuttryckte det, "Det finns en betydande överlappning mellan underrättelsenivåerav de smartaste björnar och de dummaste turister. "
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Kycklingen som clucks högljudda är det som mest sannolikt att visa uppvid ånga montörer "picknick.
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Kon är ingenting annat än en maskin som gör gräs passar för oss människor att äta.
		-- John McNulty

%
Daily PlanetSUPERMAN SPARAR dessert!Planer på att "äta det senare"
		-- John McNulty

%
Den tidiga fågeln får kaffet kvar från kvällen innan.
		-- John McNulty

%
Historien om varje större Galactic Civilization tenderar att passera igenomtre distinkta och igenkännbara faser, de Survival, undersökning ochFörfining, annars känd som hur, varför, och var faser. FörExempelvis är den första fasen kännetecknas av frågan "Hur kan vi äta?"den andra med "Varför äter vi?" och den tredje med "Var ska vi äta lunch?".
		-- Hitchhiker's Guide to the Galaxy

%
Kosher Dill uppfanns 1723 av Joe Kosher och Sam dill. Det ärden enskilt mest populära pickle variation i dag, hade hela den friavärld av man, kvinna och barn lika. En häpnadsväckande 350 miljarder kosherdill äts varje år, i genomsnitt ut till nästan 1/4 pickle per personper dag. New York Times matkritikern Mimi Sheraton säger "Den kosher dillverkligen förändrat mitt liv. Jag brukade få äta McDonalds hamburgare ochdricka Iron City Lite, och sedan jag stötte på den kosher dill pickle.Jag insåg att det fanns mycket mer att haute cuisine skulle jag någonsin trott.Och nu, bara titta på mig. "
		-- Hitchhiker's Guide to the Galaxy

%
De män satt läppja deras te i tystnad. Efter en stund klutz sade,"Livet är som en skål med gräddfil.""Som en skål med gräddfil?" frågade den andra. "Varför?""Hur ska jag veta det? Är jag en filosof?"
		-- Hitchhiker's Guide to the Galaxy

%
Den mest utsökta topp i matkultur erövras när du gör rätt genom enskinka, en skinka, i själva karaktären av bearbetning som skett sedan den senasteDet gick på egna ben, kombinerar i sin smak dofter av rökig höstskogen, moderns mjukhet jordnära fält som levereras av sina grödor barn,den wineyness en sen sol, den intima kyss gödsling regn, ochbita av brand. Du måste skiva den tunt, nästan lika tunn som denna sida hålleri dina händer. Tillverkningen av en skinka middag, som skapandet av en gentleman,börjar en lång, lång tid före evenemanget.från "Kongressen eate It Up"
		-- W. B. Courtney, "Reflections of Maryland Country Ham",

%
Den mest anmärkningsvärda om min mamma är att under trettio år hon tjänstgjordefamiljen bara resterna. Den ursprungliga måltiden har aldrig påträffats.
		-- Calvin Trillin

%
"The National Association of Theater Koncessionshavare rapporterade att i1986 var 60% av alla godis som säljs i biografer såldes till Roger Ebert. "
		-- D. Letterman

%
Antalet fötter i en gård är direkt proportionell mot den framgångav grillen.
		-- D. Letterman

%
Antalet lakrits gumballs du få ut av en gumball maskinökar i direkt proportion till hur mycket du hatar lakrits.
		-- D. Letterman

%
Det enda som är bättre än kärlek är mjölk.
		-- D. Letterman

%
Anledningen till att det kallas "Grape Nötter" är att det innehåller "dextros", som äribland även kallad "druvsocker", och även på grund av "Grape Nötter" ärcatchier, när det gäller marknadsföring, än "en korsning mellan Gerbil Mat ochGrus ", vilket är vad det smakar.
		-- Dave Barry, "Tips for Writer's"

%
Scenen: i en stor, målad öken, står inför en cowboy hans häst.Cowboy: "Ja, du har varit en ganska bra hoss, antar jag Hardworkin"..Inte den snabbaste nötkreatur jag någonsin kommer acrost, men ... "Häst: "Nej, dum, inte foder * tillbaka * Jag sa att jag ville ha en matnings * påse *..
		-- Dave Barry, "Tips for Writer's"

%
Problemet med att äta italiensk mat är att fem eller sex dagar senaredu är hungrig igen.
		-- George Miller

%
Vägen till en mans mage är genom hans matstrupe.
		-- George Miller

%
Det finns tre möjliga delar till ett datum, varav minst två skall varaerbjuds: underhållning, mat och kärlek. Det är brukligt att börja enserie av datum med en hel del underhållning, en måttlig mängdmat, och ett blott antydan om kärlek. Som mängden ömhetökar, underhållning kan minskas proportionellt. närtillgivenhet är underhållning, vi inte längre kalla det dating. Under ingaomständigheter kan maten utelämnas.
		-- Miss Manners' Guide to Excruciatingly Correct Behaviour

%
Det finns tillfällen när sanningen är konstigare än fiktion och lunch tid är enav dem.
		-- Miss Manners' Guide to Excruciatingly Correct Behaviour

%
Det finns tjugofem personer kvar i världen, och tjugosju avdem är hamburgare.
		-- Ed Sanders

%
Det finns mer enkelhet i den man som äter kaviar på impuls än iman som äter Grape-Nuts på principen.
		-- G. K. Chesterton

%
Det finns ingen sincerer kärlek än kärleken till mat.
		-- George Bernard Shaw

%
Det finns alltid gratis ost i en råttfälla.
		-- George Bernard Shaw

%
Det finns inget som ansiktet av ett barn att äta en Hershey bar.
		-- George Bernard Shaw

%
Tretton vid ett bord är otur endast när värdinnan har endast tolv kotletter.
		-- Groucho Marx

%
Detta är Betty Frenel. Jag vet inte vem du ska ringa men jag kan inte nå minMat-a-holics partner. Jag är på Vido är på min andra pizza med korvoch svamp. Jim, komma och hämta mig!
		-- Groucho Marx

%
Detta är National Non-Dairy Creamer veckan.
		-- Groucho Marx

%
... Denna strävan efter excellens sträcker sig in i människors personligalever också. När 80-talet människor köper något, köper de den bästa, sombestäms av (1) pris och (2) bristande tillgänglighet. Eighties folk köperimporterade tandtråd. De köper gourmet bakpulver. Om en 80-pargår till en restaurang där de har gjort en reservation tre veckor iavancera, och de informeras om att deras bord är tillgänglig, de förföljaomedelbart, det är inte en utmärkt restaurang eftersom de vet. Omdet var, det skulle ha en enorm skara Excellence inriktade personersom de själva väntar deras personsökare går ut som syrsor inatt. En utmärkt restaurang skulle inte ha en tabell redo omedelbartför någon under rangen av Liza Minnelli.
		-- Dave Barry, "In Search of Excellence"

%
Gå ner i vikt, äta mindre; att gå upp i vikt, äta mer; om du baravill behålla, gör vad du gjorde.Bronx kost är en legitim system för livsmedelsbehandling visar attMat ska användas en krycka och vilken mat kan vara den mest effektiva ifrämja andlig och känslomässig tillfredsställelse. För första gången, eneater kunde omedelbart förstå sambandet mellan lindra depression ochMallomars, och förstå varför en älskare gräl är inte så illa om det finns enpint glass i närheten.
		-- Richard Smith, "The Bronx Diet"

%
Att se slaktaren slap biff, innan han lade den på blocket,och ge sin kniv en skärpning, var att glömma frukost direkt. Det varangenäm, också - det var verkligen - att se honom skära bort det, så slät och saftig.Det fanns ingenting vilde på bar gärning, även om kniven var stor och angelägen;det var ett konstverk, hög konst; Det var delikatess av beröring, klarhetton, skicklig hantering av ämnet, fina skuggning. Det var triumftänka över materien; ganska.
		-- Dickens, "Martin Chuzzlewit"

%
Tom hungriga, tid att äta lunch.
		-- Dickens, "Martin Chuzzlewit"

%
För sentEtt stort antal turkies [sic] gick till San Francisco igår medde två klockan båtar. Om deras avsikt med att gå ner var att delta iThanksgiving festligheter i den staden, skulle de anländer "dagen efteraffären ", och naturligtvis tyvärr besviken därigenom.
		-- Sacramento Daily Union, November 29, 1861

%
Två jordnötter gick genom New York. Man blev överfallen.
		-- Sacramento Daily Union, November 29, 1861

%
Grönsaker är vad mat äter.Frukt är grönsaker som lura dig genom att smaka bra.Fisk är snabbrörliga grönsaker.Svampar är vad som växer på grönsaker när maten är klar med dem.
		-- Meat Eater's Credo, according to Jim Williams

%
Vegetarianer varning! Du är vad du äter.
		-- Meat Eater's Credo, according to Jim Williams

%
Servitör: "Te eller kaffe, mina herrar?"1 kund: "I have te."2nd kund: "Jag också - och vara säker på att glaset är rent!"(Servitör utgångar, returer)Servitör: ". Två te Vilken bad om rent glas?"
		-- Meat Eater's Credo, according to Jim Williams

%
Vakna upp och lukta på kaffet.
		-- Ann Landers

%
Vilka matar dessa munsbitar vara!
		-- Ann Landers

%
Vad är mat till en, är att andra bitter gift.
		-- Titus Lucretius Carus

%
Vad som är viktigt är mat, pengar och möjligheter för att ha dödat av sinfiender. Ge en man dessa tre saker och du kommer inte att höra mycket squawkingav honom.
		-- Brian O'Nolan, "The Best of Myles"

%
När en person går på en diet, är det första han förlorar sitt humör.
		-- Brian O'Nolan, "The Best of Myles"

%
När allt annat misslyckas, ÄTA !!!
		-- Brian O'Nolan, "The Best of Myles"

%
När min hjärna börjar rulla från mina litterära arbeten, jag gör en tillfälligost dopp.
		-- Ignatius Reilly

%
"När du vaknar på morgonen, Puh", sa Nasse äntligen"Vad är det första du säger till dig själv?""Vad blir det till frukost?" sa Puh. "Vad säger du, Nasse?""Jag säger, jag undrar vad som kommer att hända spännande idag?" sa Nasse.Puh nickade eftertänksamt. "Det är samma sak", sade han.
		-- Ignatius Reilly

%
När du äta ute och du misstänker att något är fel, är du förmodligen rätt.
		-- Ignatius Reilly

%
Vart går du för att få anorexi?
		-- Shelley Winters

%
Även om det kan vara sant att en bevakad pott aldrig kokar, det du intehålla ett öga på kan göra en förskräcklig röra av kaminen.
		-- Edward Stevenson

%
Den som berättar en lögn inte kan vara renhjärtade - och endast de renhjärtadekan göra en god soppa.
		-- Ludwig Van Beethoven

%
Varför så många livsmedel kommer förpackade i plast? Det är ganska kuslig.
		-- Ludwig Van Beethoven

%
Varför de kallar en snabb en snabb, när det går så långsamt?
		-- Ludwig Van Beethoven

%
Utan kaffe han inte kunde arbeta, eller åtminstone han inte kunde har arbetat isätt han gjorde. Förutom papper och pennor, tog han med sig överallt som enoumbärlig artikel av utrustning kaffemaskinen, som var mindreviktigare för honom än hans bord eller sin vita dräkt.
		-- Stefan Zweigs, Biography of Balzac

%
Utan glass liv och berömmelse är meningslösa.
		-- Stefan Zweigs, Biography of Balzac

%
Du kan alltid säga julen är här när du börjar fåotroligt tät, aluminiumfolie-och-Band- inslagna klumpar i posten. fruitcakesgöra perfekta presenter eftersom Postal Service har inte kunnat hitta ett sätt attskada dem. De evigt, till stor del eftersom ingen någonsin äter dem. IFaktum är att många smarta människor rädda fruitcakes de får och skicka dem tillbakade ursprungliga givare nästa år; vissa fruitcakes har gått tillbakaoch tillbaka i hundratals år.Det enklaste sättet att göra en fruktkaka är att köpa en mörkare kaka, sedan pundnågra gamla, hård frukt i den med en klubba. Var noga med att bära skyddsglasögon.
		-- Dave Barry, "Simple, Homespun Gifts"

%
Du behöver inte sy med en gaffel, så jag ser ingen anledning att äta med stickor.
		-- Miss Piggy, on eating Chinese Food

%
Du första föräldrar av den mänskliga rasen ... som förstört dig för ett äpple,Vad skulle du ha gjort för en truffled kalkon?
		-- Brillat-savarin, "Physiologie du Gout"

%
Du vet att du har en liten lägenhet när Rice Krispies eko.
		-- S. Rickly Christian

%
Du vet att du är en lite fett om du har bristningar på din bil.
		-- Cyrus, Chicago Reader 1/22/82

%
Du måste äta i vår cafeteria. Du kan äta smuts billig där !!!!
		-- Cyrus, Chicago Reader 1/22/82

%
Du bör tips servitören $ 10, minus $ 2 om han talar om sitt namn, en annan $ 2om han hävdar att det kommer att vara hans nöje att hjälpa dig och en annan $ 2 för varje"Special" han beskriver som involverar förvirrande begrepp som "schalottenlök," och $ 4Om menyn innehåller ordet "fixin s." I många restauranger, innebär detta attservitör kommer faktiskt skyldig dig pengar. Om du reser med ett barn i åldernsex månader till tre år, bör du lämna ett ytterligare belopp som är lika medtvå gånger räkningen för att kompensera för det faktum att de måste tabankett ut och bränna den, eftersom sprickorna är inklämt fast med gobbetstillverkad av delvis tuggade tidigare restaurang rullar mättade med baby spotta.I New York, tips taxi föraren $ 40 om han inte nämna hans hemorrojder.
		-- Dave Barry, "The Stuff of Etiquette"

%
Ditt sinne är den del av dig som säger,"Why'n'tcha äta det piece of cake?"... Och sedan, tjugo minuter senare, säger"Du vet, om jag var du, jag skulle inte ha gjort det!"
		-- Steven and Ondrea Levine

%
