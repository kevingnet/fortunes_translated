En burk sparris, 73 duvor, några LIVE ammunition och en frusen daquiri !!
		-- Bob Violence

%
En dvärg passerar ut någonstans i Detroit!
		-- Bob Violence

%
En välväxt KATOLSK SCHOOL är nervösa i min dräkt ..
		-- Bob Violence

%
Ett storögt, oskyldig UNICORN, redo fint på en äng fylldmed syrener, klubbor och små barn på HUSH av skymning ??
		-- Bob Violence

%
Egentligen, vad jag skulle vilja är en liten leksak rymdskepp !!
		-- Bob Violence

%
Allt jag kan tänka på är en platta av organiska PRUNE chips tramparav en armé av svartmuskiga, italienska LOUNGE SINGERS ...
		-- Bob Violence

%
Helt plötsligt, jag vill kasta över min lovande agerar karriär, växaen lång svart skägg och bära en baseballhatten !! ... Även om jag vet inte varför !!
		-- Bob Violence

%
Allt liv är en Blur av republikaner och kött!
		-- Bob Violence

%
Okej, urartar dig! Jag vill ha det här stället evakueras på 20 sekunder!
		-- Bob Violence

%
Under hela denna tid har jag tittar på en RYSKA MIDGET sodomize en huskatt!
		-- Bob Violence

%
Okej, du !! Imitera en WOUNDED SEAL pleading efter en parkeringsplats !!
		-- Bob Violence

%
Jag tillsammans med en förälder eller vårdnadshavare?
		-- Bob Violence

%
Jag valde ännu?
		-- Bob Violence

%
Är jag i forskarskolan ännu?
		-- Bob Violence

%
Jag snatteri?
		-- Bob Violence

%
Amerika!! Jag såg allt !! Kräkningar! Vinka! JERRY FALWELLING indin void rör av UHF glömska !! SAFEWAY i sinnet ...
		-- Bob Violence

%
En luft pommes frites genomsyrar mina näsborrar !!
		-- Bob Violence

%
En bläck-LING? Visst - TA en !! Köpte du varje kommunist UNIFORMER ??
		-- Bob Violence

%
En italiensk kammar sitt hår i en förort DES MOINES!
		-- Bob Violence

%
Och dessutom är min bowling genomsnitt oklanderlig !!!
		-- Bob Violence

%
ANN JILLIAN HÅR gör LONI Andersons hår ser ut som RICARDOMontalbán HÅR!
		-- Bob Violence

%
Är den ångade PLOMMON fortfarande i hårtorken?
		-- Bob Violence

%
Är vi lever eller på bandet?
		-- Bob Violence

%
Är vi på STRIKE ännu?
		-- Bob Violence

%
Är vi där än?
		-- Bob Violence

%
Är vi där än? Mitt sinne är en ubåt !!
		-- Bob Violence

%
Är du mentalt här på Pizza Hut ??
		-- Bob Violence

%
Säljer du NYLON oljekällor ?? Om så är fallet, kan vi använda två dussin !!
		-- Bob Violence

%
Är du fortfarande en alkoholist?
		-- Bob Violence

%
Som president Jag måste gå dammsuga min myntsamling!
		-- Bob Violence

%
Awright, som en av er gömde min penisavund?
		-- Bob Violence

%
Barbara Stanwyck gör mig nervös !!
		-- Bob Violence

%
Barbie säger Ta Quaaludes i gin och gå till ett diskotek direkt!Men Ken säger Woo-woo !! Ingen kredit på "Mr Liquor" !!
		-- Bob Violence

%
BARRY ... Det var den mest hjärtevärmande återgivande av "Jag gjorde det MINSÄTT "jag någonsin hört !!
		-- Bob Violence

%
Som en skallig hjälte är nästan lika FESTLIGT som TATUERAD knockwurst.
		-- Bob Violence

%
Bela Lugosi är mitt co-pilot- ...
		-- Bob Violence

%
BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI-BI
		-- Bob Violence

%
... Bleakness ... ödeläggelse ... plast gafflar ...
		-- Bob Violence

%
Bo Derek förstört mitt liv!
		-- Bob Violence

%
Pojke, är jag glad att det är bara 1971 ...
		-- Bob Violence

%
Pojkar, har du alla valts ut att lämna th "PLANET i 15 minuter !!
		-- Bob Violence

%
Men de gick till MARS runt 1953 !!
		-- Bob Violence

%
Men var han mogen nog kväll på lesbisk maskerad?
		-- Bob Violence

%
Kan jag har en impuls objekt i stället?
		-- Bob Violence

%
Kan du skicka en bönor kaka?
		-- Bob Violence

%
Ketchup och senap överallt! Det är den mänskliga Hamburger!
		-- Bob Violence

%
Chubby Checker hade bara en kyckling smörgås i centrala DULUTH!
		-- Bob Violence

%
Civilisationen är kul! Hur som helst, det håller mig upptagen !!
		-- Bob Violence

%
Rensa tvättomat !! Denna virvel-o-matic hade bara en härdsmälta !!
		-- Bob Violence

%
Koncentrera dig på th'cute, Li'l TECKNAD killar! Kom ihåg SERIALTAL!! Följ Whipple AVE. UTGÅNG!! Har en gratis PEPSI !! SvängVÄNSTER på th'HOLIDAY INN !! GÅ kredit världen !! GÖR MIG ETT ERBJUDANDE !!!
		-- Bob Violence

%
GRATTIS! Nu ska jag göra tunt beslöjade kommentarer omVÄRDIGHET, självkänsla och finna SANN FUN i höger kammare ??
		-- Bob Violence

%
Innehåll: 80% polyester, 20% DACRONi ... servitrisen uniform skjulTANDSTEN sås som en 8 "med 10" GLANSIG ...
		-- Bob Violence

%
Kan jag ha en överdos?
		-- Bob Violence

%
Har en italiensk kranförare uppleva bara ohämmade känsla ien MALIBU badtunna?
		-- Bob Violence

%
Gjorde jag en FEL sak ??
		-- Bob Violence

%
Sa jag att jag var en sardin? Eller en buss ???
		-- Bob Violence

%
Har jag sälja ut ännu ??
		-- Bob Violence

%
Hittade du en DIGITAL titta på i ditt låda velveeta?
		-- Bob Violence

%
Har du flyttar en hel del KOREAN stek knivar denna resa, Dingy?
		-- Bob Violence

%
DIDI ... är att en marsian namn, eller är vi i ISRAEL?
		-- Bob Violence

%
Gjorde jag inte köpa en 1951 Packard från dig sista mars i Kairo?
		-- Bob Violence

%
Disco olja Bussing kommer att skapa en bultande naugahide rörledning rinnandedirekt till tropikerna från mattan producerande regioner och devalvera dollarn!
		-- Bob Violence

%
Har jag en livsstil än?
		-- Bob Violence

%
Vet ni vi just passerat igenom ett svart hål i rymden?
		-- Bob Violence

%
Har du exakt vad jag vill ha i en pläd poindexter bar bat ??
		-- Bob Violence

%
Vill du "ANBUDS vittles"?
		-- Bob Violence

%
Tror du att "Monkees" ska få gas på udda eller jämna dagar?
		-- Bob Violence

%
Har någon från Peoria har en kortare uppmärksam än mig?
		-- Bob Violence

%
gör din omklädningsrum har tillräckligt SPARRIS?
		-- Bob Violence

%
INTE gå !! Jag är inte Howard Cosell !! Jag vet polska skämt ... VÄNTA !!Gå inte !! JAG ÄR Howard Cosell! ... Och jag vet inte polska skämt !!
		-- Bob Violence

%
Inte slog mig !! Jag är i Twilight Zone !!!
		-- Bob Violence

%
Inte SANFORISERA mig !!
		-- Bob Violence

%
Oroa dig inte, ingen verkligen lyssnar på föreläsningar i Moskva, antingen! ...FRANSKA, historia, ADVANCED Analys, programmering, SVARTSTUDIER, sociobiology! ... Finns det några frågor ??
		-- Bob Violence

%
Edwin Meese gjorde mig bära CORDOVANS !!
		-- Bob Violence

%
Eisenhower !! Din MIMEOGRAFERA ​​maskin upsets min mage !!
		-- Bob Violence

%
Antingen BEKÄNNA nu eller vi gå till "folkets domstol" !!
		-- Bob Violence

%
Alla får fri BORSCHT!
		-- Bob Violence

%
Alla kommer någonstans !! Det är förmodligen en loppmarknad eller enkatastrof film !!
		-- Bob Violence

%
Överallt ser jag jag ser negativitet och ASFALT ...
		-- Bob Violence

%
Ursäkta mig, men det gjorde jag inte berätta det finns inget hopp för överlevnadOFFSET PRINTING?
		-- Bob Violence

%
Känslor är överlappande över mig !!!
		-- Bob Violence

%
Slutligen, Zippy kör sin 1958 RAMBLER METROPOLITAN i fakultetenmatsal.
		-- Bob Violence

%
Först ska jag ge dig alla svar på dagens test ... Såbara att koppla in din SONY Walkman och slappna av !!
		-- Bob Violence

%
LURAS dig! Absorbera EGO shattering impuls strålar, polyester poltroon !!
		-- Bob Violence

%
för konstgjorda smakämnen !!
		-- Bob Violence

%
Fyra tusen olika magnater, puckelpist & NABOBS är skuttade i mittgotisk solarium !!
		-- Bob Violence

%
FRYST FÖRRÄTTER kan slungas av medlemmar av motsatta SWANSON Sects ...
		-- Bob Violence

%
FUN aldrig behöva säga att du är SUSHI !!
		-- Bob Violence

%
Gee, jag känner typ av ljus i huvudet nu, vet jag kan inte göra minparabolantenn betalningar!
		-- Bob Violence

%
Gibble, kluckande, vi accepterar DIG ...
		-- Bob Violence

%
Ge dem radarstyrda SKEE-ball körfält och velveeta BURRITOS !!
		-- Bob Violence

%
Gå på, Emote! Jag växte upp på tanke ballonger !!
		-- Bob Violence

%
God natt, alla ... Nu måste jag gå administrera FÖRSTA HJÄLPEN minsällskapsdjur Leisure Suit !!
		-- Bob Violence

%
Hårvatten, vänligen !!
		-- Bob Violence

%
En halv sinne är en fruktansvärd sak att avfall!
		-- Bob Violence

%
Ge mig ett par skinnbyxor och en CASIO tangentbord - Jag lever för idag!
		-- Bob Violence

%
Har alla fick halvah spridda över sina vrister ?? ... Nu är dettid till "HA EN NAGEELA" !!
		-- Bob Violence

%
... Han dominerar den dekadenta SUBWAY scenen.
		-- Bob Violence

%
Han är MELBA-VARA ... ängeln tårta ... XEROX honom ... XEROX honom -
		-- Bob Violence

%
Han förmodligen bara vill ta över mina celler och sedan EXPLODERA inuti migsom ett fat rinnande hackad lever! Eller kanske han villPSYCHOLIGICALLY Derbes mig tills jag har inget att invända mot en högerMilitära maktövertagandet av min lägenhet !! Jag antar att jag borde ringa Al Pacino!
		-- Bob Violence

%
HELLO KITTY gäng terroriserar staden, familj stickered till döden!
		-- Bob Violence

%
Hej, alla, jag är en människa !!
		-- Bob Violence

%
Hej, GORRY-O !! Jag är ett geni från Harvard !!
		-- Bob Violence

%
Hallå. Jag vet att skilsmässor bland ogifta katolska Alaskan honor !!
		-- Bob Violence

%
Hallå. Bara gå längs och försöker att inte tänka på dina tarmarär nästan fyrtio GÅRDAR LONG !!
		-- Bob Violence

%
Hej ... järnridå? Skicka över en korv pizza! World War III? Nej tack!
		-- Bob Violence

%
Hallå? Lavemang Bondage? Jag ringer för att jag vill vara lycklig, antar jag ...
		-- Bob Violence

%
Här är jag på loppis men ingen köper mina urinprov flaskor ...
		-- Bob Violence

%
Här är jag i 53 f Kr och allt jag vill är en dill pickle !!
		-- Bob Violence

%
Här är jag i bakre LUKT- lobule men jag kan inte se CARL SAGANnågonstans!!
		-- Bob Violence

%
Här är vi i Amerika ... när vi samla arbetslöshet?
		-- Bob Violence

%
Vänta en minut !! Jag vill ha en skilsmässa !! ... Du inte Clint Eastwood !!
		-- Bob Violence

%
Hej, servitör! Jag vill ha en ny skjorta och en hästsvans med citron sås!
		-- Bob Violence

%
Hiccuping och darrande i soptippar i New Jersey som någraberusade Kål lappar DOLL, hosta i linje vid FIORUCCI'S !!
		-- Bob Violence

%
Hmmm ... en lamslagen REVISOR med en falafel smörgås träffas av enTråd CAR ...
		-- Bob Violence

%
Hmmm ... En hash-sångare och en skelögd kille sover på en ödeö, när ...
		-- Bob Violence

%
Hmmm ... ett knappnålshuvud, under en jordbävning, stöter på ett ALL-MIDGETFIDDLE ORCHESTRA ... ha ... ha ...
		-- Bob Violence

%
Hmmm ... en arrogant bukett med en subtil antydan av POLYVINYLKLORID ...
		-- Bob Violence

%
Håll MAYO och passera COSMIC MEDVETENHET ...
		-- Bob Violence

%
Hurra, Ronald !! Nu kan du gifta dig med Linda Ronstadt också !!
		-- Bob Violence

%
Hur får jag hem?
		-- Bob Violence

%
Hur förklarar du Wayne Newton makt över miljontals? Det är th "MOUSTACHE... Har du någonsin märkt th "sätt utstrålar UPPRIKTIGHET, ärlighet & VÄRME?Det är en mustasch dig vill ta hem och presentera för Nancy Sinatra!
		-- Bob Violence

%
Hur många retured murare från FLORIDA är ute köper RITABrynen just nu ??
		-- Bob Violence

%
Hur går det i dessa MODULAR LOVE ENHETER ??
		-- Bob Violence

%
Hur är frun? Är hon hemma njuter kapitalismen?
		-- Bob Violence

%
hubub, hubub, hubub, hubub, hubub, hubub, hubub, hubub, hubub, hubub.
		-- Bob Violence

%
HUGH BEAUMONT dog 1982 !!
		-- Bob Violence

%
MÄNSKLIGA repliker är insatt i kar av näringsmässiga jäst ...
		-- Bob Violence

%
Jag har alltid kul eftersom jag ut ur mitt sinne !!!
		-- Bob Violence

%
Jag är en gelé munk. Jag är en gelé munk.
		-- Bob Violence

%
Jag är ett trafikljus, och Alan Ginzberg kidnappade min tvätt i 1927!
		-- Bob Violence

%
Jag täckt med ren vegetabilisk olja och jag skriver en bästsäljare!
		-- Bob Violence

%
Jag är djupt oroad och jag vill ha något bra för frukost!
		-- Bob Violence

%
Jag har FUN ... Jag undrar om det är NET FUN eller grov FUN?
		-- Bob Violence

%
Jag är inte en mutter ....
		-- Bob Violence

%
Jag utser dig ambassadör till Fantasy Island !!!
		-- Bob Violence

%
Jag tog min bowlingklot - och vissa läkemedel !!
		-- Bob Violence

%
Jag kan inte bestämma vilka fel väg att göra först !! Jag undrar om BOBGuccione har dessa problem!
		-- Bob Violence

%
Jag kan inte tänka på det. Det går inte med häckar i form avLITTLE LULU - eller robotar som gör BRICKS ...
		-- Bob Violence

%
Jag kräver STRAFFRIHET!
		-- Bob Violence

%
Jag beställt inte någon WOO-WOO ... Kanske YUBBA ... Men ingen WOO-WOO!
		-- Bob Violence

%
Jag tror inte att det verkligen finns en gasbrist .. Jag tror att det är allt baraen STOR HOAX på den del av plastskylt försäljare - att sälja fler nummer !!
		-- Bob Violence

%
... Jag vet inte varför, men plötsligt, jag vill diskutera sjunkande I.Q.NIVÅER med ett blått band SENAT underkommitté!
		-- Bob Violence

%
Jag vet inte varför jag sa att ... jag tror att det kom från fyllningarna imina bakre kindtänderna ...
		-- Bob Violence

%
... Jag gillar inte Frank Sinatra eller sina barn.
		-- Bob Violence

%
Jag förstår inte HUMOR av The Three Stooges !!
		-- Bob Violence

%
Jag känner ... HALSVEN ...
		-- Bob Violence

%
Jag mår bättre om världens problem nu!
		-- Bob Violence

%
Jag känner mig som en våt parkeringsautomat på Darvon!
		-- Bob Violence

%
Det känns som jag delar en `` majs DOG '' med NIKITA Khruschev ...
		-- Bob Violence

%
Det känns som jag är i en toalettskål med en häftstift i min panna !!
		-- Bob Violence

%
Jag känner delvis hydrerad!
		-- Bob Violence

%
Jag fylla mitt avfallsbehållare industri med gamla exemplar av "VAKTTORN"och sedan lägga till HAWAIIAN PUNCH till toppen ... De ser NICE på gården ...
		-- Bob Violence

%
Jag antar att det var en dröm ... eller en episod av Hawaii Five-O ...
		-- Bob Violence

%
Jag antar att ni fick stora muskler från att göra alltför mycket STUDERAR!
		-- Bob Violence

%
Jag hade ett leasingavtal på en OEDIPUS COMPLEX tillbaka i '81 ...
		-- Bob Violence

%
Jag hade pannkaka makeup för brunch!
		-- Bob Violence

%
Jag har en liten skål i mitt huvud
		-- Bob Violence

%
Jag har en mycket bra dental plan. Tack.
		-- Bob Violence

%
Jag har en vision! Det är en RANCID dubbel Fishwich på en anrikad BUN !!
		-- Bob Violence

%
Jag har accepterat Provolone i mitt liv!
		-- Bob Violence

%
Jag har många tabeller och diagram ..
		-- Bob Violence

%
... Jag har läs instruktionerna ...
		-- Bob Violence

%
- Jag har sett FUN -
		-- Bob Violence

%
Jag har sett dessa ÄGG fyllmedel i min Supermarket ... Jag har lästINSTRUKTIONER ...
		-- Bob Violence

%
Jag har befogenhet att stoppa produktionen på alla TONÅRS- SEX komedier !!
		-- Bob Violence

%
Jag måste köpa en ny "Dodge GIRIGBUK" och två dussin Jordache JEANS eftersommin viewscreen är "Ett användarvänligt" !!
		-- Bob Violence

%
Jag har inte varit gift i över sex år, men vi hade sexuell rådgivningvarje dag från Oral Roberts !!
		-- Bob Violence

%
Jag hoppas att jag köpte rätt relish ... ZZZZZZZZZ ...
		-- Bob Violence

%
Jag hoppas något gott kom med posten i dag så jag har en anledning att leva !!
		-- Bob Violence

%
Jag hoppas att `` Eurythmics "praxis preventivmedel ...
		-- Bob Violence

%
Jag hoppas att ni miljonärer har roligt! Jag investerade bara halva livbesparingar i jäst !!
		-- Bob Violence

%
Jag uppfann skydiving 1989!
		-- Bob Violence

%
Jag gick scientology på en loppmarknad !!
		-- Bob Violence

%
Jag glömde bara hela mitt livsfilosofi !!!
		-- Bob Violence

%
Jag fick bara min PRINCE bildekal ... Men nu kan jag inte minnas vem han är ...
		-- Bob Violence

%
Jag hade bara en näsoperation !!
		-- Bob Violence

%
Jag hade min hela tarmkanalen belagd med TEFLON!
		-- Bob Violence

%
Jag bara hörde sjuttiotalet var över !! Och jag var bara att få kontaktmed min Leisure Suit !!
		-- Bob Violence

%
Jag tänkte bara något om en padda!
		-- Bob Violence

%
Jag kaiser roll ?! Hur bra är en Kaiser rulle utan lite cole slawpå sidan?
		-- Bob Violence

%
Jag vet ett skämt !!
		-- Bob Violence

%
Jag vet hur man gör SPECIALEFFEKTER !!
		-- Bob Violence

%
Jag vet th'MAMBO !! Jag har en två toner CHEMISTRY UPPSÄTTNING !!
		-- Bob Violence

%
Jag vet saker om Troy Donahue som inte ens skrivas !!
		-- Bob Violence

%
Jag lämnade min plånbok i badrummet !!
		-- Bob Violence

%
Jag gillar hur ENDAST munnen flytta ... De ser ut att dö OYSTERS
		-- Bob Violence

%
Jag gillar din SNOOPY POSTER !!
		-- Bob Violence

%
- Jag älskar Katrinka eftersom hon kör en Pontiac. Vi ska bortnu. Jag matade katten.
		-- Bob Violence

%
Jag älskar Rock'n Roll! Jag memorerade alla orden till "WIPE-OUT" i1965 !!
		-- Bob Violence

%
Jag behöver diskutera återköp bestämmelser åtminstone sex studio SLEAZEBALLS !!
		-- Bob Violence

%
Jag en gång dekorerade min lägenhet helt i tio fot sallad gafflar !!
		-- Bob Violence

%
Jag äger sju åttondelar av alla artister i centrala Burbank!
		-- Bob Violence

%
Jag lägga undan min kopia av "BOWLING världen" och tänka på vapenkontrolllagstiftning...
		-- Bob Violence

%
Jag representerar en sardin !!
		-- Bob Violence

%
Jag begär en helg i Havanna med Phil Silvers!
		-- Bob Violence

%
... Jag ser toalettsitsar ...
		-- Bob Violence

%
Jag valde E5 ... men jag har inte hört "Sam Sham och Pharoahs"!
		-- Bob Violence

%
Jag luktar en RANCID corn dog!
		-- Bob Violence

%
Jag luktar som en våt minska klinik på Columbus Day!
		-- Bob Violence

%
Jag tror att jag är en overnight sensation just nu !!
		-- Bob Violence

%
... Jag tror att jag skulle bättre gå tillbaka till mitt skrivbord och leksak med några vanligaMissförstånd ...
		-- Bob Violence

%
Jag tror att jag ska döda mig genom att hoppa ut ur denna 14 STORY fönstret medanläsning Erica Jong poesi !!
		-- Bob Violence

%
Jag tror att min karriär är förstört!
		-- Bob Violence

%
Jag brukade vara en fundamentalist, men då jag hörde om HIGHStrålningsnivåer och köpte en encyklopedi !!
		-- Bob Violence

%
... Jag vill ha en COLOR T.V. och en vibrerande säng !!!
		-- Bob Violence

%
Jag vill ha en vegetariska burrito att gå ... med EXTRA MSG !!
		-- Bob Violence

%
Jag vill ha en WESSON OIL leasing !!
		-- Bob Violence

%
Jag vill ha en annan omskrivning på min ceasar sallad !!
		-- Bob Violence

%
Jag vill öron! Jag vill ha två runda svarta öron att göra mig varm 'n säker !!
		-- Bob Violence

%
... Jag vill fyrtiotvå TRYNEL FLOATATION system installerade inomSex och en halv timmar !!!
		-- Bob Violence

%
Jag vill ordförandeskapet så dåligt jag kan redan smaka smårätter.
		-- Bob Violence

%
Jag vill klä dig som Tallulah Bankhead och täcker dig med vaselinoch vete tunnar ...
		-- Bob Violence

%
Jag vill döda alla här med en gullig färgrik Vätebomb !!
		-- Bob Violence

%
... Jag vill utföra hjärnverksamhet med Tuesday Weld !!
		-- Bob Violence

%
Jag vill läsa min nya dikt om fläsk hjärnor och yttre rymden ...
		-- Bob Violence

%
Jag vill så glad, venerna i nacken STÅ UT !!
		-- Bob Violence

%
Jag vill att du ska memorera samlade dikter av Edna St. Vincent Millay... TILLBAKA !!
		-- Bob Violence

%
Jag vill att du ska organisera mina KONDITORI brickor ... mitt te-burkar är glänsande ibildning som en rad med DRUM Majorettes - vänligen inte vara rasande med mig -
		-- Bob Violence

%
Jag föddes i en Hostess Cupcake fabriken innan den sexuella revolutionen!
		-- Bob Violence

%
Jag gjorde munkar och nu är jag på en buss!
		-- Bob Violence

%
Jag önskar att jag var en sex-svalt manikyr hittades död i Bronx !!
		-- Bob Violence

%
Jag önskar att jag var på en Cincinnati gathörn håller en ren hund!
		-- Bob Violence

%
Jag undrar om jag någonsin skulle kunna komma igång i kredit världen?
		-- Bob Violence

%
Jag undrar om jag borde berätta om mitt tidigare liv som en FÄRDIGFRÄMLING?
		-- Bob Violence

%
Jag undrar om jag ska lägga mig i ESCROW !!
		-- Bob Violence

%
Jag undrar om det finns något gott i kväll?
		-- Bob Violence

%
Jag skulle vilja att urinera i en ovular, porslin pool -
		-- Bob Violence

%
Jag skulle vilja MIN databas julienned och wokade!
		-- Bob Violence

%
Jag skulle vilja ha lite SKRÄPMAT ... och då vill jag vara ensam -
		-- Bob Violence

%
Jag ska äta något som är klarblå !!
		-- Bob Violence

%
Jag ska visa er min telexnummer om du visar mig din ...
		-- Bob Violence

%
Jag är en fuschia bowlingklot någonstans i Bretagne
		-- Bob Violence

%
Jag är ett geni! Jag vill att bestrida meningsbyggnad med Susan Sontag !!
		-- Bob Violence

%
Jag är en atomubåt i polarisen och jag behöver en Kleenex!
		-- Bob Violence

%
Jag är också mot BODY surfning !!
		-- Bob Violence

%
Jag är också pre-HÄLLS pre-mediterade och prerafaelitiska !!
		-- Bob Violence

%
Jag är ANN LANDERS !! Jag kan snatta !!
		-- Bob Violence

%
Jag byta kanal ... Men allt jag får är reklam för "RONCOMIRAKEL BAMBOO hushållsprodukter "!
		-- Bob Violence

%
Jag är ständigt förvånad över th'breathtaking effekterna av vinderosion !!
		-- Bob Violence

%
Jag är definitivt inte i Omaha!
		-- Bob Violence

%
Jag FÖRTVIVLAD ... Jag hoppas att det är något friterad enligt dennaminiatyr Kupolformigt stadion ...
		-- Bob Violence

%
Jag klär i en illasittande murgröna LEAGUE PASSAR !! För sent...
		-- Bob Violence

%
Jag är EMOTIONELL nu eftersom jag har MERCHANDISING SLAG !!
		-- Bob Violence

%
Jag inkapslad i slemhinnan i en ren fläskkorv !!
		-- Bob Violence

%
Jag är glad att jag kom ihåg att XEROX alla mina undertröjor !!
		-- Bob Violence

%
Jag glider över en kärnavfalls DUMP nära Atlanta, Georgia !!
		-- Bob Violence

%
Jag har en Big Bang Theory !!
		-- Bob Violence

%
Jag har en matiné KRIS!
		-- Bob Violence

%
Jag har en religiös upplevelse ... och jag tar inte några droger
		-- Bob Violence

%
Jag har en avdragsgill upplevelse! Jag behöver en energikris !!
		-- Bob Violence

%
Jag har en känslomässig utbrott !!
		-- Bob Violence

%
Jag har en emotionellt utbrott !! Men, eh, varför finns det en våffla imin pyjamas POCKET ??
		-- Bob Violence

%
Jag har vackra tankar om fadd fruar självbelåten ochrika affärsjurister ...
		-- Bob Violence

%
Jag har kul att lifta till Cincinnati eller Far Rockaway !!
		-- Bob Violence

%
... Jag föreställa sig en sinnlig GIRAFF, cavorting i det inre rummetav en kosher Deli -
		-- Bob Violence

%
Jag är i direkt kontakt med många avancerade roliga BEGREPP.
		-- Bob Violence

%
Jag är i SOFTWARE!
		-- Bob Violence

%
Jag mediterar på formaldehyd och asbesten läcker in i minPERSONLIGT UTRYMME!!
		-- Bob Violence

%
Jag är mentalt övertrasseras! Vad är det SIGN längre fram? Var är RODSTERLING när du verkligen behöver honom?
		-- Bob Violence

%
Jag är inte en iransk !! Jag röstade för Dianne Feinstein !!
		-- Bob Violence

%
Jag är inte tillgänglig för en kommentar ..
		-- Bob Violence

%
Jag låtsas att jag drar i en öring! Gör jag det rätt ??
		-- Bob Violence

%
Jag låtsas att vi alla tittar Phil Silvers istället RicardoMontalban!
		-- Bob Violence

%
Jag tyst läsning senaste numret av "BOWLING WORLD" medan min fruoch två barn står tyst vid ...
		-- Bob Violence

%
Jag betyget PG-34 !!
		-- Bob Violence

%
Jag får ett kodat meddelande från Eubie BLAKE !!
		-- Bob Violence

%
Jag är RELIGIOUS !! Jag älskar en man med en POSTISCH !! Utrusta mig med missiler !!
		-- Bob Violence

%
Jag rapporterar för arbetsuppgift som en modern människa. Jag vill göra det latinska Hustle nu!
		-- Bob Violence

%
Jag rakar !! JAG RAKA !!
		-- Bob Violence

%
Jag sitter på min hastighet QUEEN ... För mig, det är roligt ... Jag är VARMT... Jag är VIBRATORS ...
		-- Bob Violence

%
Jag tänker om digital avläsningssystem och datorgenereradeBILDKONSTELLATIONER ...
		-- Bob Violence

%
Jag är helt FÖRTVIVLAD över situationen i Libyen och priset på kyckling ...
		-- Bob Violence

%
Jag använder min X-RAY VISION för att erhålla en sällsynt glimt av INREHur denna POTATIS !!
		-- Bob Violence

%
Jag bär PAMPERS !!
		-- Bob Violence

%
Jag är våt! Jag är vild!
		-- Bob Violence

%
Jag är ung ... jag är frisk ... jag kan vandra THRU CAPT Grogan'S ländrygg!
		-- Bob Violence

%
Jag Zippy PINHEAD och jag är helt engagerad i festläge.
		-- Bob Violence

%
Jag har en kusin som arbetar i Garment District ...
		-- Bob Violence

%
Jag har en idé!! Varför jag inte stirra på dig så hårt, du glömtPERSONNUMMER!!
		-- Bob Violence

%
Jag har läst sju miljoner böcker !!
		-- Bob Violence

%
... Ich bin in einem dusenjet ins Jahr 53 vor chr ... ich lande imAntiken Rom ... einige Gladiatoren spielen scrabble ... ich riechePIZZA ...
		-- Bob Violence

%
Om en person är känd i detta land, måste de gå på vägen förMånader åt gången och har sitt namn felstavat på sidan av enVINTHUND SCENICRUISER !!
		-- Bob Violence

%
Om vald, lovar Zippy till varje amerikansk en 55-årig houseboy ...
		-- Bob Violence

%
Om jag blir vald ingen någonsin kommer att behöva göra sin tvätt igen!
		-- Bob Violence

%
Om jag blir vald, kommer betongbarriärer runt VITA HUSET varaersättas med smakfulla skum kopior av Ann-Margret!
		-- Bob Violence

%
Om jag kände någon mer sofistikerad skulle jag dö förlägenhet!
		-- Bob Violence

%
Om jag hade en tops, kan jag förhindra th "kollaps av förhandlingar !!
		-- Bob Violence

%
... Om jag hade hjärtsvikt just nu, kan jag inte vara en mer lyckosam man !!
		-- Bob Violence

%
Om jag drar den här växeln I be Rita Hayworth !! Eller en scientolog!
		-- Bob Violence

%
om det glittrar, sluka det !!
		-- Bob Violence

%
Om vårt beteende är strikt, behöver vi inte kul!
		-- Bob Violence

%
Om Robert Di Niro mördar Walter Slezak, kommer Jodie Foster gifta Bonzo ??
		-- Bob Violence

%
År 1962 kunde man köpa ett par hajskinn BYXOR, med en "ContinentalBälte, "för $ 10,99 !!
		-- Bob Violence

%
I Newark de tvättomater är öppen 24 timmar om dygnet!
		-- Bob Violence

%
INSIDE, jag har samma personlighetsstörning som LUCY RICARDO !!
		-- Bob Violence

%
Inuti jag redan GRÅT!
		-- Bob Violence

%
Är en tatuering verklig, som en trottoarkant eller ett slagskepp? Eller är vi lider i Safeway?
		-- Bob Violence

%
Är han MAGIC INCA bär en groda på sina axlar ?? Är grodanhans Guide ?? Det är märkligt att en hund körs redan på rulltrappan ...
		-- Bob Violence

%
Är det 1974? Vad för Nattvarden? Kan jag tillbringar min college fond i envild eftermiddag ??
		-- Bob Violence

%
Är det ren i andra dimensioner?
		-- Bob Violence

%
Är det nouvelle cuisine när 3 Oliver kämpar med en pilgrimsmussla i enplatta sås MORNAY?
		-- Bob Violence

%
Är något VIOLENT kommer att hända med en soptunna?
		-- Bob Violence

%
Är detta en out-take från "BRADY GRUPPEN"?
		-- Bob Violence

%
Kommer detta att innebära RAW mänsklig extas?
		-- Bob Violence

%
Är detta TERMINAL kul?
		-- Bob Violence

%
Är detta raden för den senaste nyckfull jugoslaviska drama som ocksågör du vill gråta och ompröva Vietnamkriget?
		-- Bob Violence

%
Är inte detta mitt STOP ?!
		-- Bob Violence

%
Det betyder inte en sak om du inte har fått det SWING !!
		-- Bob Violence

%
Det var ett skämt!! Förstår?? Jag tog emot meddelanden från David Letterman !!YOW !!
		-- Bob Violence

%
Det är mycket roligt att leva ... Jag undrar om min säng görs?!?
		-- Bob Violence

%
Det är ingen användning ... Jag har gått till "CLUB MED" !!
		-- Bob Violence

%
Det är uppenbart ... pälsarna nådde aldrig ISTANBUL ... Du var en EXTRAi nyinspelningen av "TOPKAPI" ... Gå hem till din fru ... Hon görFATTIGA RIDDARE!
		-- Bob Violence

%
Det är okej - Jag är en intellektuell, alltför.
		-- Bob Violence

%
Det är sköljcykeln !! De har alla ignorerade sköljningen !!
		-- Bob Violence

%
JAPAN är en underbar planet - Jag undrar om vi någonsin kommer att nå sin nivåav jämförande shopping ...
		-- Bob Violence

%
Jesuitpräster dejta diplomatiska tjänstemän !!
		-- Bob Violence

%
Jesus är min POSTMÄSTARE GENERAL ...
		-- Bob Violence

%
Ungar, inte brutto mig ... "Adventures med mental hygien" kan varatransporteras för långt!
		-- Bob Violence

%
Ungar, sju baslivsmedel grupper är GUM, PUFF bakverk, pizza,Pesticider, antibiotika, Nutra-Sweet och MJÖLKblindgångare !!
		-- Bob Violence

%
Tvätt är den femte dimensionen !! ... Um ... um ... e 'tvättmaskinär ett svart hål och rosa strumpor är bussförare som bara blev !!
		-- Bob Violence

%
LBJ, LBJ, hur många skämt sa du idag ??!
		-- Bob Violence

%
Leona, jag vill erkänna saker till dig ... jag vill WRAP dig i en rödROBE trimmas med POLYVINYL KLORID ... Jag vill tömma ASKKOPPAR ...
		-- Bob Violence

%
Låt mig göra min tribute till nätstrumpor ...
		-- Bob Violence

%
Låt oss alla visa mänsklig omsorg om Reverand månens juridiska svårigheter !!
		-- Bob Violence

%
Låt oss skicka ryssarna defekta livsstil tillbehör!
		-- Bob Violence

%
Livet är en popularitetstävling! Jag är UPPFRISKANDE CANDID !!
		-- Bob Violence

%
Som jag alltid säger - ingenting kan slå bratwurst här i Düsseldorf !!
		-- Bob Violence

%
Loni Anderson hår bör legaliseras !!
		-- Bob Violence

%
Titta djupt in i öppningarna !! Ser du några älvor eller EDSELS ... eller enGROGG?? ...
		-- Bob Violence

%
Titta in i mina ögon och försöka glömma att du har en Macys betalkort!
		-- Bob Violence

%
Se! En stege! Kanske det leder till himlen, eller en smörgås!
		-- Bob Violence

%
SE!! Tystlåten amerikanska tonåringar bär MADRAS shorts och "Flock avSeagulls "frisyrer!
		-- Bob Violence

%
Gör mig att se ut som Linda Ronstadt igen !!
		-- Bob Violence

%
Mary Tyler Moores SJUNDE MAKA bär min DACRON linne i enbilliga hotell i Honolulu!
		-- Bob Violence

%
Kanske kan vi måla Goldie Hawn en rik berlinerblått -
		-- Bob Violence

%
Meryl Streep är min förlossningsläkare!
		-- Bob Violence

%
MMM-MM !! Så detta är BIO-NEBULATION!
		-- Bob Violence

%
Mmmmmm-MMMMMM !! En platta med ångande bitar av en PIG blandas med denstrimlor av FLERA KYCKLINGAR !! ... Oh Jösses!! Jag är på väg att svälja enAvrivna delen av en COW vänstra ben indränkt i bomullsfröolja ochSOCKER!! ... Låt oss se ... Nästa, I have grunden och upp kött av söta,Baby lamm stekta i de smälta, fettvävnad från ett varmblodigtdjur någon gång petted !! ... YUM !! Det var bra!! Till efterrätt,Jag har en tofu burgare med Bean GRODDAR på en sten marken, HELAVETE BUN !!
		-- Bob Violence

%
Herr och fru PED, kan jag låna 26,7% av rayon textilproduktion avden indonesiska övärlden?
		-- Bob Violence

%
Min moster MAUREEN var en militär rådgivare till Ike & Tina Turner !!
		-- Bob Violence

%
Min biologiska VÄCKARKLOCKA bara gick ... Det har ljudlös DOZEFUNKTION och komplett kök !!
		-- Bob Violence

%
Min Code of Ethics är semestrar på berömda Schroon Lake i upstate New York !!
		-- Bob Violence

%
Mina öron är borta !!
		-- Bob Violence

%
Mitt ansikte är nytt, min licens har gått ut, och jag är under en läkares vård !!!!
		-- Bob Violence

%
Min frisyr är helt traditionella!
		-- Bob Violence

%
Min inkomst är alla engångs!
		-- Bob Violence

%
Min LESLIE GORE rekord är trasig ...
		-- Bob Violence

%
Mitt liv är en uteplats roligt!
		-- Bob Violence

%
Mitt sinne är en potatisåker ...
		-- Bob Violence

%
Mitt sinne gör askkoppar i Dayton ...
		-- Bob Violence

%
Min näsa känns som en dålig Ronald Reagan film ...
		-- Bob Violence

%
Min näsa är stel!
		-- Bob Violence

%
... Mina byxor bara gick på en vild framfart genom en Long Island Bowling Alley !!
		-- Bob Violence

%
Mina byxor bara gick i gymnasiet i Carlsbad Caverns !!!
		-- Bob Violence

%
Min polyvinyl cowboy plånbok gjordes i Hongkong av Montgomery Clift!
		-- Bob Violence

%
Min morbror Murray erövrade Egypten 53 f Kr Och jag kan bevisa det också !!
		-- Bob Violence

%
Min vaselin körs ...
		-- Bob Violence

%
NANCY !! Varför är allt RED ?!
		-- Bob Violence

%
NATHAN ... dina föräldrar var i en CARCRASH !! De ogiltigförklaras - deKollapsade De hade inga SÅGAR ... De hade inga pengar maskiner ... Degjorde piller i TORFTIG gräs kjolar ... Nathan, jag emuleras dem ... mende var OFF-KEY ...
		-- Bob Violence

%
NEWARK har rezoned !! DES MOINES har rezoned !!
		-- Bob Violence

%
Bröstvårtor, gropar, knogar, Nickles, rynkor, finnar !!
		-- Bob Violence

%
Inte SENSUOUS ... bara "SPRALLIG" ... och i behov av tandvård ... smärta !!!
		-- Bob Violence

%
Nu är jag deprimerad ...
		-- Bob Violence

%
Nu tror jag att jag nådde bara tillståndet av högt blodtryck som kommer JUSTInnan du ser TOTAL på Safeway kassadisken!
		-- Bob Violence

%
Nu förstår jag innebörden av "Gänget"!
		-- Bob Violence

%
Nu Jag blir ofrivilligt blandas närmare CLAM DIP medBROKEN plast gafflar i det !!
		-- Bob Violence

%
Jag är nu att koncentrera sig på en specifik tank strid mot slutet av andra världskriget!
		-- Bob Violence

%
Nu jag har fadd tankar om den vackra, runda fruarHollywoodfilm Moguls inneslutna i plexiglas CARS och att närma sigav småpojkar som säljer frukt ...
		-- Bob Violence

%
Nu KEN och BARBIE är permanent ADDICTED till sinnesförändrande droger ...
		-- Bob Violence

%
Nu är mina känslomässiga resurser är starkt åtagit sig att 23% av smältningoch raffineringsindustrin i delstaten Nevada !!
		-- Bob Violence

%
Nu när jag har min "äpple", jag förstår COST REDOVISNING !!
		-- Bob Violence

%
Nu ska vi SKICKA UT för QUICHE !!
		-- Bob Violence

%
Naturligtvis, du förstå om plädar i centrifugeringen -
		-- Bob Violence

%
Herregud - SUN bara föll i Yankee Stadium !!
		-- Bob Violence

%
Oh jag fattar!! "Stranden går på", va, SONNY ??
		-- Bob Violence

%
Okej ... Jag kommer hem för att skriva "JAG HATAR Rubiks kub HANDBOK FÖRDöd katt älskare "...
		-- Bob Violence

%
OKEJ!! Slå på ljudet endast för TRYNEL mattor, fullt utrustatR.V.'S och FLOATATION SYSTEMS !!
		-- Bob Violence

%
Allsidiga MEDVETENHET ?? Åh Yeh !! Först behöver fyra liter JELL-Ooch en stor NYCKEL !! ... Jag tror att du tappar th'WRENCH i JELL-O som omDet var en smak, eller en ingrediens ... ... eller ... Jag ... um ... VAR ÄRtvättmaskiner?
		-- Bob Violence

%
Vid närmare eftertanke kanske jag ska värma upp några bakade bönor och titta på RegisPhilbin ... Det är fantastiskt att vara vid liv !!
		-- Bob Violence

%
Å andra sidan, kan livet vara en ändlös parad av transsexuellQuiltning BIN ombord på ett kryssningsfartyg till Disneyworld om vi bara låter det !!
		-- Bob Violence

%
På vägen är ZIPPY ett knappnålshuvud utan ett syfte, men aldrig utan en punkt.
		-- Bob Violence

%
En gång i tiden, fyra AMFIBISK HOG ringer attackerade en familj avFörsvarslös, KÄNSLIGA myntsamlare och fällde sin egendomVÄRDEN !!
		-- Bob Violence

%
En gång, det var inte roligt ... Det var innan menyplanering, FASHIONuttalanden eller NAUTILUS utrustning ... Då, 1985 ... FUN varhelt kodad i denna lilla MICROCHIP ... Det innehåller 14.768 vagtroliga sitcom-piloter !! Vi var tvungna att vänta fyra miljarder år, men viäntligen Jerry Lewis, MTV och ett stort urval av creme-fylldasnacktårtor!
		-- Bob Violence

%
En Fishwich kommer upp !!
		-- Bob Violence

%
Ett liv att leva för alla mina barn i en annan värld alla dagar av våra liv.
		-- Bob Violence

%
ONE: Jag kommer att donera min hela "BABY HUEY" serietidning samling tillcentrala PLASMA CENTER ...TVÅ: Jag kommer inte att starta ett band som heter "khadafy & THE HIT SQUAD" ...TRE: Jag kommer aldrig torktumling min foxterrier igen !!
		-- Bob Violence

%
... Eller var du kör PONTIAC som tutade på mig i MIAMI förra tisdag?
		-- Bob Violence

%
Fader vår som är i himmelen ... Jag ber uppriktigt att någon på dettaTabellen kommer att betala för min strimlad VAD och engelska muffins ... och ävenlämna ett generöst tips ....
		-- Bob Violence

%
över i västra Philadelphia en valp kräkningar ...
		-- Bob Violence

%
OVER underpass! Under överfart! Runt framtiden och inte kan repareras !!
		-- Bob Violence

%
Ursäkta mig, jag talar engelska?
		-- Bob Violence

%
Ursäkta mig, men vet du vad det innebär att vara verkligen en med din monter!
		-- Bob Violence

%
Peggy Fleming stjäl BASKET bollar att mata barn i Vermont.
		-- Bob Violence

%
Människor förödmjuka en salami!
		-- Bob Violence

%
PIZZA!!
		-- Bob Violence

%
Placera mig på en bufferträknare när du förringa flera bellhops iTrianon Room !! Låt mig en av dina DOTTERBOLAG!
		-- Bob Violence

%
Kom hem med mig ... Jag har Tylenol !!
		-- Bob Violence

%
Psyko ?? Jag trodde att detta var en naken rap session !!!
		-- Bob Violence

%
Punk rock !! Disco duck !! PREVENTIVMEDEL!!
		-- Bob Violence

%
Snabb, sjunga mig BUDAPEST NATIONAL ANTHEM !!
		-- Bob Violence

%
SLÄKT!!
		-- Bob Violence

%
Kom ihåg att i 2039, kommer MOUSSE och pasta vara tillgängliga endast av recept !!
		-- Bob Violence

%
Rhapsody in lim!
		-- Bob Violence

%
SANTA CLAUS kommer ner en brandstege bära ljusa blå benvärmare... Han scrubs påven med en mild tvål eller rengöringsmedel i 15 minuter,starring Jane Fonda !!
		-- Bob Violence

%
Skicka dina frågor till `` ASK ZIPPY '', Box 40474, San Francisco, Kalifornien94140, USA
		-- Bob Violence

%
SHHHH !! Jag hör SIX Tatuerade truckförare gungade motorblock itomma oljefat ...
		-- Bob Violence

%
Ska jag göra mitt BOBBIE VINTON medley?
		-- Bob Violence

%
Ska jag få låst i PRINCICAL'S OFFICE idag - eller har en vasektomi ??
		-- Bob Violence

%
Ska jag börja med den tid jag bytte personligheter med en BEATNIKfrisör eller min underlåtenhet att hänvisa fem tonåringar att en bra OKULIST?
		-- Bob Violence

%
Skriv i min framställning.
		-- Bob Violence

%
Så det här är hur det känns att vara potatissallad
		-- Bob Violence

%
Så, om vi omvandlar utbudssidan soja FUTURES i högavkastande T-BILLINDIKATORER, kommer PRE-inflationsriskerna krympa till en hastighet av 2Shoppingrundor per AUBERGINE !!
		-- Bob Violence

%
Någon i Dayton, Ohio är sälja begagnade mattor till en serbokroatiska
		-- Bob Violence

%
Någon gång under 1993 Nancy Sinatra kommer att leda en oblodig kupp på Guam !!
		-- Bob Violence

%
Någonstans i centrala BURBANK en prostituerad är kokning en LAMB CHOP !!
		-- Bob Violence

%
Någonstans i en förort till Honolulu, har en arbetslös piccolo piska upp ensats av illegal psilocybin chop suey !!
		-- Bob Violence

%
Någonstans i Tenafly, New Jersey, är en kiropraktor tittar "Låt denBeaver "!
		-- Bob Violence

%
Sprida jordnötssmör påminner mig om opera !! Jag undrar varför?
		-- Bob Violence

%
Tailfins !! ... klick ...
		-- Bob Violence

%
Talar Pinhead Blues:Åh, förlorade jag min `` HELLO KITTY '' DOLL och jag får dålig mottagning på kanal    Tjugosex !!Th'HOSTESS Fabriken closin "ner och jag bara hört Zasu Pitts har varit    Död sedan många år .. (sniff)Min PLATTFORM skokollektion var tuggas upp av th "hund, Alexander Haig    kommer inte att låta mig ta en dusch "til påsk ... (snurf)Så jag gick till köket, men WALNUT PANELING whup mig upp mah HAID !!    (På nej, nej, nej .. Heh, heh)
		-- Bob Violence

%
TAPPNING? Du POLITIKER! Inser ni inte att slutet av "WashCykel "är en värdefull ögonblick för de flesta människor ?!
		-- Bob Violence

%
Tex SEX! HOME hjul! Det droppar av kaffe !! Ta mig tillMinnesota men inte genera mig !!
		-- Bob Violence

%
Th MIND är Pizza Palace of th "SOUL
		-- Bob Violence

%
Tack Gud!! ... Det är HENNY Youngman !!
		-- Bob Violence

%
Uppskattning av den genomsnittliga visuella graphisticator enbart är värthela suaveness och dekadens som vimlar !!
		-- Bob Violence

%
Hela den kinesiska kvinnor volleybollag alla delar en personlighet -och har sedan födseln !!
		-- Bob Violence

%
Det faktum att 47 personer är skriker och svetten forsande ner minRyggraden tämligen angenäm !!
		-- Bob Violence

%
Falafel SANDWICH landar på mitt huvud och jag bli vegetarian ...
		-- Bob Violence

%
... Motorvägen är gjord av kalk JELLO och min HONDA är en barbequeuedOSTRON! Yum!
		-- Bob Violence

%
Koreakriget måste ha varit kul.
		-- Bob Violence

%
... De Mysterians är här med min CORDUROY SOAP skålen !!
		-- Bob Violence

%
Osmonds! Ni är alla Osmonds !! Att kasta upp på en motorväg i gryningen !!!
		-- Bob Violence

%
Pillsbury Doughboy gråter till ett slut på Burt Reynolds filmer !!
		-- Bob Violence

%
Den rosa strumpor var ursprungligen från 1952 !! Men de gick till MARSomkring 1953 !!
		-- Bob Violence

%
Samma WAVE håller kommer in och kollapsar som en rayon MUU-MUU ...
		-- Bob Violence

%
Det finns ingen sanning. Det finns ingen verklighet. Finns det ingen konsekvens.Det finns inga absoluta uttalanden. Jag är mycket sannolikt fel.
		-- Bob Violence

%
Det finns en liten bild av ED MCMAHON gör dåliga saker att Joan Riversi en $ 200.000 MALIBU BEACH HOUSE !!
		-- Bob Violence

%
Det finns tillräckligt med pengar för att köpa 5000 burkar Noodle-Roni!
		-- Bob Violence

%
"Det är mörka tider för alla mänsklighetens högsta värdena!""Dessa är mörka tider för frihet och välstånd!""Det är bra tider att sätta dina pengar på skurk att sparka CRAPut ur Megaton MAN! "
		-- Bob Violence

%
Dessa konserver vara tvångsmatas till Pentagon !!
		-- Bob Violence

%
De kollapsade ... som nunnor på gatan ... de hade ingen tonåringöverklagande!
		-- Bob Violence

%
Detta KÖNLÖS PIG egentligen handlar mitt blod ... Han är så ... så ... BRÅDSKANDE !!
		-- Bob Violence

%
"Detta är ett jobb för BOB VÅLD och avskum, den otroligt korkat MUTANT HUND."
		-- Bob Violence

%
Detta är en utan krusiduller flyg - håll th "Canadian bacon !!
		-- Bob Violence

%
Detta måste vara en bra fest - bröstkorgen är smärtsamt trycks uppmot någons MARTINI !!
		-- Bob Violence

%
... Det måste vara hur det är att vara en högskoleexamen !!
		-- Bob Violence

%
Denna pizza symboliserar hela min EMOTIONELL ÅTERHÄMTNING !!
		-- Bob Violence

%
Detta PORCUPINE vet hans ZIPCODE ... Och han har "VISA" !!
		-- Bob Violence

%
Detta toppar av min partygoing upplevelse! Någon som jag inte gillar ärprata med mig om en värmande europeisk film ...
		-- Bob Violence

%
De är inte Winos - det är min jonglör, mitt aerialist, mitt svärdSwallower, och min LATEX NOVELTY LEVERANTÖR !!
		-- Bob Violence

%
Tusentals dagar civila ... har producerat en ... känsla förestetiska moduler -
		-- Bob Violence

%
Idag, tre Winos från DETROIT sålde mig ett inramat foto av TAB HUNTERinnan hans makeover!
		-- Bob Violence

%
Tår, knän, bröstvårtor. Tår, knän, bröstvårtor, KNOGAR ...Bröstvårtor, gropar, knogar, Nickles, rynkor, finnar !!
		-- Bob Violence

%
Tony Randall! Är ditt liv en uteplats på FUN ??
		-- Bob Violence

%
Uh-oh - varför jag plötsligt att tänka på en ärevördig religiös ledareplaskar på en FORTLAUDERDALE helgen?
		-- Bob Violence

%
Hoppsan!! Jag glömde att underkasta sig OBLIGATORISK urinanalys!
		-- Bob Violence

%
HOPPSAN!! Jag satte på "STORA rakt på tågkollisioner av 50-talet" avmisstag!!!
		-- Bob Violence

%
HOPPSAN!! Jag tror KEN är ÖVER DUE på hans R.V. BETALNINGAR och han har enNERVOUS FÖRDELNING också !! Haha.
		-- Bob Violence

%
Hoppsan!! Jag har för mycket roligt !!
		-- Bob Violence

%
HOPPSAN!! Vi är av bildelar och gummivaror!
		-- Bob Violence

%
Begagnade häftklamrar är bra med soja!
		-- Bob Violence

%
Vicariously uppleva några anledning att leva !!
		-- Bob Violence

%
Rösta för mig - jag är väl avsmalnande, halv-spänd, ogenomtänkta och uppskjuten skatt!
		-- Bob Violence

%
Vänta ... Detta är en rolig sak eller slutet av livet i Petticoat Junction ??
		-- Bob Violence

%
Var min SOY SLÄNTRAR utelämnats i th'RAIN? Det smakar riktigt bra !!
		-- Bob Violence

%
Vi är nu njuter total ömsesidig samverkan i en imaginär barrel ...
		-- Bob Violence

%
Vi har olika mängder hår -
		-- Bob Violence

%
Vi gick bara det civila hår patrull!
		-- Bob Violence

%
Vi lägger två kopior av tidningen People i en mörk, fuktig husbil.45 minuter senare Cyndi Lauper framträder bär en fågelbur på huvudet!
		-- Bob Violence

%
Tja, här är jag i Amerika .. Jag gillar det. Jag hatar det. Jag gillar det. jagHatar det. Jag gillar det. Jag hatar det. Jag gillar det. Jag hatar det. JAG GILLAR ...Känslor sveper över mig !!
		-- Bob Violence

%
Tja, jag är en klassisk ANAL MOTTAGLIG !! Och jag letar efter ett sätt attVicariously uppleva några anledning att leva !!
		-- Bob Violence

%
Tja, jag är osynlig igen ... Jag kan lika gärna besöka LadiesRUM ...
		-- Bob Violence

%
Okej då. Jag kompromissa med mina principer på grund existentiell FÖRTVIVLAN!
		-- Bob Violence

%
Var dessa palsternacka RÄTT marinerad i tacosås?
		-- Bob Violence

%
Vilket sammanträffande! Jag är en auktoriserad "snoots av stjärnorna" dealer !!
		-- Bob Violence

%
Hur bra är en papp resväska ÄNDÅ?
		-- Bob Violence

%
Vad jag behöver är en mogen relation med en diskett ...
		-- Bob Violence

%
Vad jag vill veta är - papegojor vet mycket om Astro-Turf?
		-- Bob Violence

%
Vilket program de tittar på?
		-- Bob Violence

%
Vad universum är detta, vänligen ??
		-- Bob Violence

%
Vad är det för fel Sid? ... Är din dryck otillfredsställande?
		-- Bob Violence

%
När jag träffade th'POPE tillbaka i '58, skrubbade jag honom med en mild tvål ellerRENGÖRINGSMEDEL under 15 minuter. Han tycktes njuta av det ...
		-- Bob Violence

%
När denna belastning KLAR Jag tror jag ska tvätta den igen ...
		-- Bob Violence

%
När du får din Ph.D. kommer du att få möjlighet att arbeta på Burger King?
		-- Bob Violence

%
När du sa "skogrika" det påminde mig om en förfallen RENGÖRINGBILL ... Ser du inte? O'Grogan svalde en värdefulla Coin COLLECTIONoch var tvungen att mörda den ende som visste !!
		-- Bob Violence

%
Var kommer dina strumpor gå när du förlorar dem i th "WASHER?
		-- Bob Violence

%
Vart tar det vägen när du spola?
		-- Bob Violence

%
Var Sandy Duncan?
		-- Bob Violence

%
Var är th "Daffy Duck EXHIBIT ??
		-- Bob Violence

%
Var är Coke maskin? Berätta ett skämt för mig!!
		-- Bob Violence

%
Medan min HJÄRNSKÅL är nekas service i Burger King, Jesuitpräster dating diplomatiska tjänstemän !!
		-- Bob Violence

%
Medan du tuggar, tror Steven Spielbergs bankkonto ... hanskommer att ha samma effekt som två "stärkelse blockerare"!
		-- Bob Violence

%
WHO ser en BEACH KANIN snyftande på en SHAG RUG ?!
		-- Bob Violence

%
OJ!! Ken och Barbie är med för mycket roligt !! Det måste varaNegativa joner !!
		-- Bob Violence

%
Varför är dessa sportsko försäljare efter mig ??
		-- Bob Violence

%
Varför inte du någonsin in några tävlingar, Marvin ?? Vet du inte dinegen ZIPCODE?
		-- Bob Violence

%
Varför är allt gjort av Lycra Spandex?
		-- Bob Violence

%
Varför är det så att när du dör, du kan inte ta din hemmabioCENTER med dig ??
		-- Bob Violence

%
Kommer det att förbättra min KASSAFLÖDE?
		-- Bob Violence

%
Kommer det tredje världskriget hålla "famn Buddies" från luften?
		-- Bob Violence

%
Kommer detta aldrig sinande rad njutbara HÄNDELSER upphör aldrig?
		-- Bob Violence

%
Med dig kan jag vara mig själv ... Vi behöver inte Dan Rather ...
		-- Bob Violence

%
World War III? Nej tack!
		-- Bob Violence

%
Tredje världskriget kan undvikas genom att ansluta sig till en strikt klädkod!
		-- Bob Violence

%
Wow! Se!! En herrelös köttbulle !! Låt oss intervjua det!
		-- Bob Violence

%
Xerox din lunch och lämna in den under "sexualbrottslingar"!
		-- Bob Violence

%
Ja, men jag ser påskharen i skintight läder på en IRONMAIDEN konsert?
		-- Bob Violence

%
Du kan inte skada mig !! Jag har en assumable INTECKNAR !!
		-- Bob Violence

%
Du menar nu kan jag skjuta dig i ryggen och ytterligare BLUR th "åtskillnad mellan fantasi och verklighet?
		-- Bob Violence

%
Du menar att du inte vill titta på BROTTNING från Atlanta?
		-- Bob Violence

%
Du valde Karl Malden näsa !!
		-- Bob Violence

%
Du bör alla hoppa upp och ner i två timmar medan jag besluta om en ny karriär !!
		-- Bob Violence

%
Du var s'posed att skratta!
		-- Bob Violence

%
DU!! Ge mig den sötaste, mest rosa, mest charmiga lilla VICTORIANDOCKHUS hittar du !! En gör det SNAPPY !!
		-- Bob Violence

%
Dina kinder sitta som tvilling NEKTARINER över en mun som inte känner några gränser -
		-- Bob Violence

%
Dagens ungdom! Gå med mig i ett massmöte för traditionell mentalattityder!
		-- Bob Violence

%
Yow!
		-- Bob Violence

%
Yow! Jag har roligt ännu?
		-- Bob Violence

%
Yow! Är jag i Milwaukee?
		-- Bob Violence

%
Yow! Och då kunde vi sitta på huvarna av bilar vid stoppljusen!
		-- Bob Violence

%
Yow! Är vi laid back ännu?
		-- Bob Violence

%
Yow! Är vi våt ännu?
		-- Bob Violence

%
Yow! Är du själv stekning president?
		-- Bob Violence

%
Yow! Har något dåligt händer eller är jag i en drive-in film ??
		-- Bob Violence

%
Yow! Jag gick under fattigdomsgränsen!
		-- Bob Violence

%
Yow! Jag kastade upp på mitt fönster!
		-- Bob Violence

%
Yow! Jag vill ha min näsa i ljus!
		-- Bob Violence

%
Yow! Jag vill skicka en bronserad kronärtskocka till Nicaragua!
		-- Bob Violence

%
Yow! Jag har en quadrophonic känsla av två winos ensam i ett stålverk!
		-- Bob Violence

%
Yow! Jag inbillar en surfare van fylld med sojasås!
		-- Bob Violence

%
Yow! Är min skyddsrum termit bevis?
		-- Bob Violence

%
Yow! Är detta samlag ännu ?? Är det, va, är det ??
		-- Bob Violence

%
Yow! Det är ett hål hela vägen till centrum Burbank!
		-- Bob Violence

%
Yow! Det är en del människor inne i väggen! Detta är bättre än att torka!
		-- Bob Violence

%
Yow! Kanske jag borde ha begärt för min Neutron bomb i Paisley -
		-- Bob Violence

%
Yow! Nu får jag tänka på alla dåliga saker jag gjorde till en BOWLINGBollen när jag var i högstadiet!
		-- Bob Violence

%
Yow! Nu kan vi bli alkoholister!
		-- Bob Violence

%
Yow! Dessa människor ser ut exakt som Donnie och Marie Osmond !!
		-- Bob Violence

%
Yow! Vi kommer att en ny disco!
		-- Bob Violence

%
YOW !! Alla ur genpool!
		-- Bob Violence

%
YOW !! Jag är i en mycket smart och bedårande INSANE ASYL !!
		-- Bob Violence

%
YOW !! Nu förstår jag avancerad mikrobiologi och th "nya skattereformen lagar !!
		-- Bob Violence

%
YOW !! Landet med den stigande SONY !!
		-- Bob Violence

%
YOW !! Där framme! Det är en munk HUT !!
		-- Bob Violence

%
YOW !! Vad ska hela den mänskliga rasen DO ?? Förbruka en femtedel avCHIVAS REGAL, skidor NAKEN ner MT. EVEREST, och har en vild SEX helg!
		-- Bob Violence

%
YOW !!! Jag har kul!!!
		-- Bob Violence

%
Zippy hjärnceller ansträngande att överbrygga synapser ...
		-- Bob Violence

%
