94% av kvinnorna i Amerika är vackra och resten umgås runt här.
		-- Oscar Wilde

%
En kandidat är en man som aldrig gjort samma misstag en gång.
		-- Oscar Wilde

%
En kandidat är en självisk, förtjänar kille som har fuskat någon kvinna utav en skilsmässa.
		-- Don Quinn

%
En kandidat är en unaltared hane.
		-- Don Quinn

%
En kandidat aldrig riktigt blir över tanken att han är en sak av skönhetoch en pojke för alltid.
		-- Helen Rowland

%
En dåligt äktenskap är som en häst med ett brutet ben, kan du skjutahästen, men det inte fixa benet.
		-- Helen Rowland

%
En vacker människa är ett paradis för ögonen, helvete för själen, ochskärseld för handväskan.
		-- Helen Rowland

%
En vacker kvinna är en välsignelse från himlen, men en god cigarr är en rök.
		-- Kipling

%
En vacker kvinna är en bild som driver alla åskådarna ädelt galen.
		-- Emerson

%
En pojke kan lära mycket av en hund: lydnad, lojalitet, och viktenatt vända tre gånger innan liggande.
		-- Robert Benchley

%
En pojke får vara en man när en människa behövs.
		-- John Steinbeck

%
En Chicago försäljare var på väg att checka in en St Louis hotell när han märkteen mycket charmig kvinna stirrar beundrande på honom. Han gick fram och talademed henne i några minuter, och återvände sedan till receptionen, där de kontrollerasi som Mr och MrsEfter en mycket angenäm tre dagars vistelse, närmade sig mannen frontenskrivbord och berättade clerk han checkar ut. Inom några minuter var han handedett lagförslag för $ 2500."Det måste vara ett misstag," försäljaren sade. "Jag har varit här förbara tre dagar. ""Ja, sir" expediten svarade. "Men din fru har varit här en månadoch en halv."
		-- John Steinbeck

%
En hederskodexen: aldrig närma sig en väns flickvän eller fru med ofogsom ditt mål. Det finns alltför många kvinnor i världen för att motivera den sortensohederliga beteende. Om hon är verkligen lockande.
		-- Bruce J. Friedman, "Sex and the Lonely Guy"

%
En diplomat är man som alltid kommer ihåg en kvinna födelsedag men aldrig hennes ålder.
		-- Robert Frost

%
En diplomatisk man sa till sin hustru, "Hur du förväntar mig att minnasdin födelsedag när du aldrig se någon äldre? "
		-- Robert Frost

%
En dominerande man gifte sig med en enkel wisp av en flicka. Han kom tillbaka frånhans smekmånad en luttrad man. Han hade blivit medveten om irrbloss.
		-- Robert Frost

%
En siffra med kurvor ger alltid en hel del intressanta vinklar.
		-- Robert Frost

%
En spännande Mercedes-Benz röt upp till trottoaren där en söt ung miss stodväntar på en taxi."Hej", sade mannen vid ratten. "Jag ska väst.""Så underbart," kom den svala svar. "Ge mig tillbaka en orange."
		-- Robert Frost

%
En dåre och hans honung snart skildes.
		-- Robert Frost

%
En räv är en varg som skickar blommor.
		-- Ruth Weston

%
En gentleman är en man som inte skulle slå en kvinna med hatten på.		[ Och varför inte? För varför hon har hatten på? Ed.]
		-- Evan Esar

%
En herre slår aldrig en dam med hatten på.
		-- Fred Allen

%
En flicka och en pojke bump i varandra - säkert en olycka.En flicka och en pojke bula och näsduken droppar - säkert en annan olycka.Men när en flicka ger en pojke en död bläckfisk - * _ _ _ _ att _ _ _ hade _ _ att _ _ _ _ menar _ _ _ _ _ _ _ _ _ något *.
		-- S. Morganstern, "The Silent Gondoliers"

%
En flicka med en framtid undviker man med ett förflutet.
		-- Evan Esar, "The Humor of Humor"

%
En flickas bästa vän är hennes mutter.
		-- Dorothy Parker

%
En flicka samvete inte riktigt hålla henne från att göra något wrong--det bara håller henne från att njuta det.
		-- Dorothy Parker

%
En god människa alltid vet sina begränsningar.
		-- Harry Callahan

%
Ett bra äktenskap skulle vara mellan en blind fru och döv man.
		-- Michel de Montaigne

%
En kille måste få frisk då och då så en flicka inte förlorar hennes förtroende.
		-- Michel de Montaigne

%
En hammare missar ibland sina spår - en bukett aldrig.
		-- Michel de Montaigne

%
En man är vad som är kvar av älskare efter nerven har utvunnits.
		-- Helen Rowland

%
En kvinna är en som aldrig visar hennes underkläder oavsiktligt.
		-- Lillian Day

%
En man måste alltid komma ihåg en sak om en vacker kvinna.Någonstans är någon trött på henne.
		-- Lillian Day

%
En man minns alltid hans första kärlek med särskild ömhet, men eftersom börjar att gäng dem.
		-- Mencken

%
En man kom hem tidigt för att hitta sin hustru i armarna på sin bästa vän,som svor hur mycket de var förälskade. Att tysta rasande make,älskare föreslog, "Vänner bör inte slåss, låt oss spela gin rummy. Om jag vinner,du får en skilsmässa så jag kan gifta sig med henne. Om du vinner, jag lovar att aldrig sehenne igen. Okej?""Okej", instämde mannen. "Men hur ungefär en fjärdedel en punktpå sidan för att göra det intressant? "
		-- Mencken

%
En man kan ha två, kanske tre kärleksaffärer medan han är gift. Efteratt det är fusk.
		-- Yves Montand

%
En man ser inte bakom dörren om han har stått där själv.
		-- Du Bois

%
En man i kärlek är ofullständig tills han är gift. Då han är klar.
		-- Zsa Zsa Gabor, "Newsweek"

%
En man är redan halvvägs förälskad i någon kvinna som lyssnar på honom.
		-- Brendan Francis

%
En man är som en rostig hjul på en rostig vagn,Han sjunger sin sång som han skramlar tillsammans och sedan faller han isär.
		-- Richard Thompson

%
En människa kan vara så mycket av allt som han är ingenting av någonting.
		-- Samuel Johnson

%
En man kan ibland bli förlåten kyssen som han inte har rätt,men aldrig kyssen han har inte initiativet att hävda.
		-- Samuel Johnson

%
En man sjönk till psykiater soffa och sade: "Jag har enfruktansvärda problem, doktorn. Jag har en son vid Harvard och en annan son vidPrinceton; Jag har bara begåvad var och en av dem med en ny Ferrari; jag harhem i Beverly Hills, Palm Beach och en co-op i New York; och jag harfick en blomstrande ranch i Venezuela. Min fru är en vacker ung skådespelerskasom anser mina två älskarinnor att vara hennes bästa vänner. "Psykiatern tittade på patienten, förvirrad. "Har jag saknarnågot? Det låter för mig som du inte har några problem alls. ""Men doktorn, jag bara göra $ 175 per vecka."
		-- Samuel Johnson

%
En man tog sin hustru hjortjakt för första gången. Efter att han hade gett hennevissa grundläggande instruktioner, enades de om att separera och rendezvous senare. Innanhan lämnade, han varnade henne om hon skulle föll en hjort att vara försiktig med jägare somkan slå henne till stommen och göra anspråk på döda. Om det hände, sade hanhenne, skulle hon skjuta sin pistol tre gånger i luften och han skulle komma tillhennes stöd.Strax efter att de separerat, hörde han ett enda skott, följde snabbtav den överenskomna signalen. Kör till platsen, fann han sin hustru ståendei en liten glänta med en mycket nervös man stirrar ner hennes eldröret."Han hävdar att detta är hans", sade hon, uppenbarligen mycket upprörd."Hon kan hålla det, hon kan hålla det!" den storögda mannen svarade. "JAGbara vill få min sadel tillbaka! "
		-- Samuel Johnson

%
En man vanligtvis faller förälskad i en kvinna som frågar den typ av frågorhan kan svara.
		-- Ronald Colman

%
En man gnäll till sin vän om hur han hatade att gå hem efter ensen kortspel."Du skulle inte tro vad jag går igenom för att undvika att vakna min fru,"sade han. "För det första jag döda motorn ett kvarter från huset och kustenin i garaget. Då jag öppna dörren långsamt, ta av mig skorna, ochtå till vårt rum. Men precis som jag är på väg att glida ner i sängen, hon alltidvaknar upp och ger mig fan. ""Jag gör en stor brummande när jag går hem", hans vän svarade.	"Du gör?""Visst. Jag tuta, slå igen dörren, slå på alla lampor,stampa upp till sovrummet och ge min fru en stor puss. `Hej, Alice, säger jag.`Vad sägs om en liten smooch för din gubbe?""Och vad säger hon?" hans vän frågade i misstro."Hon säger ingenting", hans kompis svarade. "Hon låtsas alltidhon sover. "
		-- Ronald Colman

%
En man stod på knä vid en grav på en kyrkogård, gråter och ber mycket högt,"Åh why..eeeee dog du ... eeeeee, Oh Why..eeeeee,varför gjorde du Di ...... eeee "Vaktmästaren går fram, förlåter sig själv och frågar artigt,"Ursäkta mig, sir, men jag har sett dig i timmar nu,bedriver på denna grav. Du måste ha varit mycket nära den avlidne. ""Nej, jag har aldrig träffat honom. Oh varför .... eeeee gjorde du dieeeeee,varför .... eeeee gjorde dig .. ""Sir, du säger att du aldrig träffat den här personen, men du fortsätta så?Tell, jag som är begravd här? ""Min frus förste man."
		-- Ronald Colman

%
En man pratar med sin bästa vän om hans äktenskap. "Du vet," hansäger: "Jag litar verkligen min fru, och jag tror att hon har alltid varit trogenmig, men det finns * alltid * att tvivel. Det finns * alltid * det lilla tvivel. ""Ja, jag vet vad du menar," hans vän svarar."Ja, kompis, jag har att lämna på en affärsresa i helgen,och jag undrar ... ja ... du skulle titta på mitt hus medan jag är borta? jag litar påhenne, det är bara att det finns * alltid * att tvivel. "Vännen gick med på att hjälpa till och två veckor senare gav sin rapport."Jag har fått en del dåliga nyheter för dig", säger vännen. "Kvällenefter att du lämnade jag såg en underlig bil dra upp framför huset. En manfick ut ur bilen och gick i huset och hade middag med din fru.Efter middagen gick de upp och jag såg din fru kyssa honom. Då, hantog av sig skjortan och hon tog av hennes blus. Och då ljuset gickut."	"*Vad hände sen?" sade mannen, hans ögon öppna bred."Ja, jag vet inte", svarade vännen, "det var för mörkt för att se.""Fan!" röt mannen. "Du ser vad jag menar? Det finns * alltid *att tvekan! "
		-- Ronald Colman

%
En man utan en kvinna är som en staty utan duvor.
		-- Ronald Colman

%
En man insvept i sig själv gör ett mycket litet paket.
		-- Ronald Colman

%
En man mĺste veta sina begränsningar.
		-- Clint Eastwood, "Dirty Harry"

%
En blygsam kvinna, klädd i hela sin grannlåt, är den mest enorma objekteti hela skapelsen.
		-- Goldsmith

%
En mor tar tjugo år för att göra en man av hennes pojke, och en annan kvinnagör narr av honom i tjugo minuter.
		-- Frost

%
En piedestal är lika mycket ett fängelse som alla små, trånga utrymmen.
		-- Gloria Steinem

%
En vacker kvinna kan göra vad som helst; en ful kvinna måste göra allt.
		-- Gloria Steinem

%
En psykiater är en kollega som ber dig en massa dyra frågordin fru ber dig för ingenting.
		-- Joey Adams

%
En påträngande romeo frågade en vacker hiss operatör, "Gör inte alla dessastannar och startar får du ganska slitna? "" Det är inte stopp och starteratt få på mina nerver, det är de idioter. "
		-- Joey Adams

%
En riktig gentleman tar aldrig baser om han verkligen måste.
		-- Overheard in an algebra lecture.

%
En romersk skild från sin hustru, som i hög grad klandras av hans vänner, somkrävde "Var hon inte kysk? Var hon inte rättvist? Var hon inte fruktbart?"håller ut sin sko, frågade dem om det inte var ny och väl gjorts.Ändå tillade han, kan ingen av er berätta var den klämmer mig.
		-- Plutarch

%
En skotte var promenera över High Street en dag bär hans kilt.När han närmade sig långt trottoaren, märkte han två unga blondiner i en röd cabrioleteyeing honom och giggling. En av dem ropade "Hej, Scotty! Vad bärsunder kilt? "Han spatserade över till sidan av bilen och frågade: "Ach, lass, är duSURE du vill veta? "Något nervöst svarade blonda ja, gjorde honverkligen vill veta.Skotten lutade närmare och anför, "Varför lass, är ingenting som bärsunder kilt, är allt i perfekt workin 'ordning! "
		-- Plutarch

%
En skarpare perspektiv på denna fråga är särskilt viktig för feministtänkte idag, eftersom en stor tendens i feminismen har konstrueratProblemet med dominans som ett drama av kvinnlig sårbarhet offer för manligaggression. Även de mer sofistikerade feministiska tänkare ofta blygabort från analysen av underkastelse, av rädsla för att att erkänna kvinnansdeltagande i maktförhållandet, ansvaret ansvarsser ut att skifta från män till kvinnor, och den moraliska segern från kvinnormän. Mer allmänt, har detta varit en svaghet radikal politik: attidealisera de förtryckta, som om deras politik och kultur var orörd avsystemet dominans, som om människor inte delta i sin egenunderkastelse. För att minska dominans till en enkel relation doer och gjort tillär att ersätta moralisk upprördhet för analys.
		-- Jessica Benjamin, "The Bonds of Love"

%
En sociolog, en psykolog och en ingenjör diskuteradeföljder och konsekvenser av en gift man har en älskarinna. Desociologen uppfattning var att det är absolut och kategoriskt oförlåtligten gift man gå miste om band av äktenskap, och engagera sig i en sådan ödmjukoch lustfyllda sysselsättningar.Psykologen uppfattning var att även moraliskt förkastligt,om man måste ha en älskarinna för att uppnå sin fulla potential som människa,sedan - ja - han kan gå vidare och välja att ha en älskarinna, så länge hanär hänsynsfull nog att hålla detta hemligt för sin hustru.Ingenjören inflikade då: "Jag tror också att, om nödvändigt,en gift man har rätt till en älskarinna. Men jag inte se varföraffären ska döljas från hustrun. Tvärtom, om affärenär ute i det fria, sedan på fredag ​​kvällar han kan tala om sin hustru att hankommer att se hans älskarinna, berätta för sin älskarinna att han kommer att vara medhans fru, sedan gå till hans kontor och få vissa arbete! "
		-- Jessica Benjamin, "The Bonds of Love"

%
En hustru varar endast för längden på äktenskapet, men en ex-fru är där* För resten av ditt liv *.
		-- Jim Samuels

%
En kvinna kan se både moraliskt och spännande - om hon ser också ut som om detvar ganska kamp.
		-- Edna Ferber

%
En kvinna kan aldrig vara för rik eller för tunt.
		-- Edna Ferber

%
En kvinna gjorde vad en kvinna skulle det bästa sättet hon visste hur.Att göra mer var omöjligt, att göra mindre, otänkbart.
		-- Dirisha, "The Man Who Never Missed"

%
En kvinna förlfräckheten som hennes skönhet har föranlett oss att vara skyldig.
		-- LeSage

%
En kvinna har fått älska en dålig man en gång eller två gånger i sitt liv för att varatacksam för en bra.
		-- Marjorie Kinnan Rawlings

%
En kvinna är som din skugga; Följ henne, hon flyger; flyga från henne, hon följer.
		-- Chamfort

%
En kvinna kan mycket väl bilda en vänskap med en man, men för att detta ska uthärda,Det måste få hjälp av en liten fysisk motvilja.
		-- Nietzsche

%
En kvinna med generös karaktär kommer att offra sitt liv tusen gångeröver för hennes älskare, men kommer att bryta med honom för alltid över en fråga omstolthet - för öppning eller stängning av en dörr.
		-- Stendhal

%
En kvinna ska inte behöva köpa sin egen parfym.
		-- Maurine Lewis

%
En kvinna utan en man är som en fisk utan en cykel.
		-- Gloria Steinem

%
En kvinna utan en man är som en fisk utan en cykel.Därför är en man utan en kvinna som en cykel utan en fisk.
		-- Gloria Steinem

%
En kvinnas bästa skyddet är lite pengar av hennes egna.
		-- Clare Booth Luce, quoted in "The Wit of Women"

%
En kvinnas plats är i huset ... och i senaten.
		-- Clare Booth Luce, quoted in "The Wit of Women"

%
En kvinna, särskilt om hon har oturen att veta något,bör dölja det så gott hon kan.
		-- Jane Austen

%
En ung man med ett mindervärdeskomplex insisterade han var bara enliten sten på stranden. Äktenskapet rådgivare sa till honom: "Om du villspara ditt äktenskap, skulle du bättre vara en liten sten. "
		-- Jane Austen

%
En ung man och hans flickvän gick längs Main Street när hon spotteden vacker diamantring i ett smycke-skyltfönster. "Wow, jag skulle verkligen älska atthar det! "Hon forsade."Inga problem", hennes kamrat svarade kasta en tegelsten genomfönstret och ta tag i ringen.Några kvarter senare, kvinnan beundrade en fullängds sable coat. "VadJag skulle ge att äga det, "sade hon, suckande."Inga problem", sa han och kastade en tegelsten genom fönstret och ta tagkappan.Slutligen vände för hemmet, passerade de en bilfirma. "Boy, skulle jag göranågot för en av dessa Rolls-Royce ", sade hon."Jösses, baby", killen stönade, "du tror att jag gjort av tegel?"
		-- Jane Austen

%
AA AAAAAAAAAaaaaaaaaaaaaaaaccccccccckkkkkk !!!!!!!!!Du brute! Knacka innan en damer rum!
		-- Jane Austen

%
Är inte ingenting en gammal man kan göra för mig men ge mig ett meddelande från en ung man.
		-- Moms Mabley

%
Underhåll är ett system som, när två personer gör ett misstag, en av demfortsätter att betala för det.
		-- Peggy Joyce

%
Underhåll är som att köpa havre för en död häst.
		-- Arthur Baer

%
Underhåll är förbannelse skrivklasser.
		-- Norman Mailer

%
Alla arvtagerskor är vackra.
		-- John Dryden

%
Alla män är likadana, men de har olika ansikten så att du kan berättadem isär.
		-- John Dryden

%
Alla de flesta män verkligen vill i livet är en hustru, ett hus, två barn och en bil,en katt, ingen kanske en hund. Eeeh, skrapa ett av barnen och lägga till en hund.Definitivt en hund.
		-- John Dryden

%
Alla män på min personal kan skriva.
		-- Bella Abzug

%
Allt arbete och ingen lön gör en hemmafru.
		-- Bella Abzug

%
Amerikanska kulturen bygger på bilen, och någon ung man löftekommer att äga en och vill resa långa sträckor i det. Följaktligen,någon ung kvinna av aspiration bör räkna med att tillbringa större delen av hennes semesteri en bil, att tränga in okända hörn. Hon behöver inte veta huratt köra men hon kommer säkert att förväntas läsa färdplanen medan hennesman kör, och om hon inte kan, eller om hon är onormalt långsam i att ge honomhjälp, hon skyldig att orsaka problem. Därför skulle du tror att högskolorsom utbildar de ljusa unga kvinnor som ska gifta sig med den ljusa ungamän som kommer att äga Cadillacs som ryta fram och tillbaka över dettakontinent skulle lära flickorna att läsa kartor. Ingen gör. De lär hundraandra värdelösa saker, men aldrig ett ord om det som kommer att orsakastörst friktion.
		-- James Michener, "Space"

%
En pilot förlovade sig två mycket vackra kvinnor på sammatid. En namngavs Edith; den andra namngivna Kate. De träffades, upptäckte dehade samma fästmö, och berättade för honom. "Ut ur våra liv du rackare. Vi skalär dig att du inte kan ha din Kate och Edith också. "
		-- James Michener, "Space"

%
En optimist är en man som ser fram emot äktenskap.En pessimist är en gift optimist.
		-- James Michener, "Space"

%
"Och vad gör ni tror att du gör ?!" röt mannen, som han kompå sin fru i sängen med en annan man. Hustrun vände sig om och log mot henneföljeslagare."Se?" Hon sa. "Jag sa ju att han var dum!"
		-- James Michener, "Space"

%
Och ändå jag borde ha dyrt gillade, jag äger, att ha rört hennes läppar; tillhar ifrågasatt henne, att hon skulle ha öppnat dem; att ha sett påfransarna hennes nedslagna ögon och aldrig tagit upp en rodnad; att ha låtitlös vågor av hår, skulle en tum av vilken vara en minnessak bortom pris:kort sagt, skulle jag ha velat, jag erkänner, att ha haft den lättastelicens av ett barn, och ändå varit man nog att känna sitt värde.
		-- Charles Dickens

%
Någon flicka kan vara glamorös; Allt du behöver göra är att stå stilla och ser dum.
		-- Hedy Lamarr

%
Varje kvinna är en volym om man vet hur man läser henne.
		-- Hedy Lamarr

%
Den som säger att han kan se genom kvinnor saknas en hel del.
		-- Groucho Marx

%
"Något annat, sir?" frågade uppmärksam piccolo försöker sitt bästaatt göra dam och herre bekväm i sin takvåning iposh hotell."Nej, tack", svarade mannen."Allt för din fru, sir?" piccolo frågade."Varför, ja, ung man," sade mannen. "Vill du ge mig envykort?"
		-- Groucho Marx

%
Som fäder går vanligen är det sällan en olycka att vara fader; ochmed tanke på den allmänna körningen söner, som sällan en olycka att vara barnlös.Det enda solid och varaktig fred mellan en man och hans hustru är, utan tvekan,en separation.
		-- Lord Chesterfield, letter to his son, 1763

%
På frågan om hur hon kände att den första kvinnan att göra en stor-league lag, honsa, "Som en gris i lera" eller ord om detta, och sedan vände ochsläppt en skvätt tobak saft från tuss av rom indränkt plugg i sinhögra kinden. Hon tuggade en sällsynt märke av plugg som kallas Stuff Det, som honlärt sig att tugga när hon spelade nicaraguanska sommar boll. Hon berättadeförfattare: "De var så betyder för mig där nere kan du inte skriva det i dintidning. Jag tog en pistol överallt jag gick, även till sängs. * Särskilt * tillsäng. Killarna var efter mig som om du inte kan tro. Det var då jag börjadetuggtobak - det spelar ingen roll hur dåligt någon behandlar dig, är det intelika dålig som detta. Detta är den värsta tugga i världen. Efter det här,allt annat är persikor och grädde. "Författarna valde Gentleman Jim,Sparrow har P.R. kille, att bita av en bit och berätta för dem hur det smakade,och där han satt och tuggade det tårarna rann ner sina gamla solbrända kinder och hankunde inte prata en stund. Sedan viskade han, "Du har tugga detta förtvå år? Gud, jag hade ingen aning om det var så svårt att vara en kvinna. "
		-- Garrison Keillor

%
Äntligen har jag hittat flickan i mina drömmar. I går kväll sade hon till mig,"Än en gång, konstigt, och den här gången * jag * vara Donnie och * du * vara Marie.
		-- Strange de Jim

%
Ungkarlar fruar och gamla pigor "barn är alltid perfekt.
		-- Nicolas Chamfort

%
I grund och botten min fru var omogen. Jag skulle vara hemma i badkaret och hon skullekomma in och sjunka mina båtar.
		-- Woody Allen

%
Var försiktig i dina förbindelser med kvinnor. Det är bättre att se påoperan med en man än i massa med en kvinna.
		-- De Maintenon

%
Vara beredda att acceptera uppoffringar. Vestal oskulder är inte så illa.
		-- De Maintenon

%
Beauty rekommenderar sällan en kvinna till en annan.
		-- De Maintenon

%
Skönhet, hjärnor, tillgänglighet, personlighet; plocka några två.
		-- De Maintenon

%
Före äktenskapet de tre små ord är "Jag älskar dig" efter äktenskapetde är "Låt oss äta ut."
		-- De Maintenon

%
Bakom varje framgångsrik man hittar en kvinna med något att bära.
		-- De Maintenon

%
Uppmanas solicitously om tillståndet i hennes hälsa blev besvärtill den gravida kvinnan vid cocktailparty. Och ännu en annan gäst gick överoch frågade, "Nå, hur mår du nuförtiden?""Inte så bra", säger den blivande modern. "Du vet, jag har missatsju eller åtta perioder nu och det börjar oroa mig. "
		-- De Maintenon

%
Ägs av någon brukade kallas slaveri - nu heter engagemang.
		-- De Maintenon

%
Benny Hill: Vill du ha en jordnöt?Girl: Nej tack, jag vill inte vara skyldig.Benny Hill: Du kommer inte att vara skyldig till en jordnöt.Det är inte som om det vore en chokladkaka eller något.
		-- De Maintenon

%
Bigami är att ha en make för många. Monogamy är densamma.
		-- De Maintenon

%
Fåglar och bin har så mycket att göra med livets fakta som svartnightgowns göra med att hålla varmt.
		-- Hester Mundis, "Powermom"

%
Pojkar är utanför intervallet någon är säker förståelse, åtminstonenär de är i åldrarna 18 månader och 90 år.
		-- James Thurber

%
Pojkar är pojkar, och så kommer en hel del medelålders män.
		-- Kin Hubbard

%
Banditer kommer att kräva dina pengar eller ditt liv, men en kvinna kommer att kräva både.
		-- Samuel Butler

%
Med alla medel gifta: Om du får en bra hustru, blir du glad; om dufå dåligt, blir du en filosof.
		-- Socrates

%
Ändra män / fruar är bara att byta problem.
		-- Kathleen Norris

%
Välj i äktenskapet bara en kvinna som du skulle välja som en vän om honvar en man.
		-- Joubert

%
Uppvaktning till äktenskap, som en mycket kvick prolog till en mycket tråkig spel.
		-- William Congreve

%
Darling: den populär form av adress som används i tala till en medlem avmotsatt kön vars namn du kan inte just nu komma ihåg.
		-- Oliver Herford

%
Kära fröken Manners:Jag bär en stor svart paraply, även om det finns bara en trettio procents chansregn. Får jag fråga en ung dam som är en främling för mig att dela sitt skydd?I morse var jag väntar på en buss i jämförande komfort, mitt paraplyskydda mig från skyfall, och märkte en attraktiv ung kvinna att fåuppblött. Jag har ofta sett henne på min busshållplats, även om vi aldrig har talat,och jag vet inte ens hennes namn. Kan jag har bett henne att komma under minparaply utan att verka kränkande?Gentle läsare:Säkert. Hänsyn till de mindre lyckligt lottade än du är alltid korrekt,även om det skulle vara mer övertygande om du slutade Joller om hurattraktiv hon är. För att inte ge bra Samaritanism ett dåligt rykte, frökenManners ber dig att låta henne två eller tre regniga dagar unmolested skyddinnan din attack.
		-- Oliver Herford

%
Kära fröken Manners:Vänligen lista några taktfull sätt att ta bort en mans saliv från ansiktet.Gentle läsare:Vänligen lista några anständiga sätt att förvärva en mans saliv i ansiktet. Omherrn sprutade du oavsiktligt att följa entusiastiskadiskurs, kan du steg tillbaka två steg, ta fram näsduken ochgå igenom motioner för att torka näsan, medan efterföljande duken tillsammansansiktet för att plocka upp vad behöver sög längs vägen. Om emellertidämnet förvärvades som ett resultat av entusiasm av en mer intimnatur, kan du försiktigt hämta det med en snärt med din rosa tunga.
		-- Oliver Herford

%
Låt inte en kvinna att be om förlåtelse, för det är bara den förstasteg. Den andra är motiverat av sig själv genom att anklagelser om dig.
		-- DeGourmont

%
Tycker du att din mamma och jag har levt bekvämt så längetillsammans om allt vi hade varit gift?
		-- DeGourmont

%
Förutsätt inte att varje ledsen ögon kvinna har älskat och förlorat - hon fårhar fått honom.
		-- DeGourmont

%
Vet inte vilken tid jag kommer tillbaka, mamma. Förmodligen snart efter att hon kastar ut mig.
		-- DeGourmont

%
Inte gifta för pengarna; du kan låna den billigare.
		-- Scottish Proverb

%
Dull kvinnor har immaculate hem.
		-- Scottish Proverb

%
Under ett besök i Amerika, var Winston Churchill inbjudna till en buffélunch där kall stekt kyckling serverades. Återvänder för en andrahjälpa, frågade han artigt, "Får jag lite bröst?""Mr Churchill", svarade värdinnan, "i det här landet vi ber omvitt kött eller mörkt kött. "Churchill ursäktade ymnigt.Följande morgon fick, damen en magnifik orkidé frånhennes hedersgäst. Den medföljande kortet läser: "Jag skulle vara mest tacksam omdu vill fästa detta på vitt kött. "
		-- Scottish Proverb

%
Ekonomer försöker fortfarande att räkna ut varför flickorna med minstprincip dra störst intresse.
		-- Scottish Proverb

%
Åttio procent av gifta män fuska i Amerika. Resten fuska i Europa.
		-- Jackie Mason

%
... Åttio år senare kunde han fortfarande minns med den unge pang av hansursprungliga glädje hans kär i Ada.
		-- Nabokov

%
Jämlikhet är inte när en kvinnlig Einstein blir befordrad till biträdandeprofessor; jämlikhet är när en kvinnlig KLANTSKALLE går framåt så snabbt som enmanlig KLANTSKALLE.
		-- Ewald Nyquist

%
Eugene d'Albert, en känd tysk kompositör, var gift sex gånger.Vid en kvällsmottagning som han deltog med sin femte hustru kortefter deras bröllop, presenterade han damen till en vän som sade artigt,"Grattis, herr d'Albert, du har sällan introducerade mig till såcharmiga hustru. "
		-- Ewald Nyquist

%
"Även i dag en man kan inte stiga upp och döda en kvinna utan känslabara lite unchivalrous ... "
		-- Robert Benchley

%
Varje människa som är högt upp gillar att tro att han har gjort det allt själv,och hustrun ler och låter det gå på det.
		-- Barrie

%
Alla ges samma mängd hormoner, vid födseln, ochOm du vill använda din för växande hår, det är bra med mig.
		-- Barrie

%
Jordbrukare i undersökningen rankade maskinhaverier Iowa State merstressande än skilsmässa.
		-- Wall Street Journal

%
Feminister vill bara mänskligheten att vara en slips.
		-- Wall Street Journal

%
Första kärleken är bara lite oförstånd och en hel del av nyfikenhet, ingen riktigtsjälvrespekt kvinna skulle dra nytta av det.
		-- George Bernard Shaw, "John Bull's Other Island"

%
Flirta är den milda konsten att göra en människa känner sig nöjd med sig själv.
		-- Helen Rowland

%
För en ung man, ännu inte: en gammal man, aldrig alls.När ska man gifta sig? En ung man, ännu inte; en äldre man, inte alls.
		-- Sir Francis Bacon, "Of Marriage and Single Life"

%
För en ung man, ännu inte: en gammal man, aldrig alls.När ska man gifta sig? En ung man, ännu inte; en äldre man, inte alls.
		-- Sir Francis Bacon, "Of Marriage and Single Life"

%
För jag svor jag skulle stanna ett år ifrån henne; ut och tyvärr!men med avbrott på dagen jag gick att göra bön.
		-- Paulus Silentiarius, c. 540 A.D.

%
För trettio år gick en man att spendera varje kväll med Mme. ___.När hans fru dog hans vänner trodde att han skulle gifta sig med henne, och uppmanadehonom att göra det. "Nej, nej", sade han: "om jag gjorde, var ska jag måstebringa min kvällar? "
		-- Chamfort

%
Fortunate är han för vilka belle mödor.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 14Låga Slag:Låt oss säga att en man och en kvinna tittar på en boxningsmatch på TV. Enav boxarna avverkas av en lågt slag. Kvinnan säger "Oh, jösses. Det måsteont. "Mannen fördubblar över och faktiskt känner smärta.Klä upp sig:En kvinna klär upp sig för att gå och handla, vattna blommorna, tömmaskräp, svara i telefonen, läsa en bok, hämta posten. En man klär uppför: bröllop, begravningar. På tal om bröllop, när reminiscing ombröllop, kvinnor talar om "ceremoni". Män skrattar om "kandidatpart".David Letterman:Män tror David Letterman är den roligaste mannen i ansiktet avJord. Kvinnor tycker att han är en genomsnittlig, halv töntigt kille som alltid har en dålig frisyr.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 16förhållanden:Först av allt, en man inte kalla en relation en relation - hanhänvisar till det som "den tid när jag och Suzie gjorde det på en semi-regulargrund".När ett förhållande tar slut, kommer en kvinna gråta och häll hennes hjärta ut tillhennes väninnor, och hon kommer att skriva en dikt med titeln "Alla Män är idioter". Sedanhon kommer att gå vidare med sitt liv.En man har lite mer problem att släppa taget. Sex månader efter det attupplösning, vid 03:00 på en lördag kväll, kommer han ringa och säga, "jag baraville låta du vet att du har förstört mitt liv, och jag kommer aldrig att förlåta dig, och jaghata dig, och du är en total floozy. Men jag vill att du ska veta att det finnsalltid en chans för oss ". Detta är känt som" Jag hatar dig / Jag älskar dig "berusad telefonsamtal, att 99% om alla män har gjort åtminstone en gång. Det finnscommunity college som erbjuder kurser för att hjälpa män komma över detta behov; tyvärr,dessa klasser sällan visa sig vara effektivt.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 17Skor:Den genomsnittliga människan har 4 par skor: löparskor, finskor,stövlar och tofflor. Den genomsnittliga kvinnan har skor 4 lager tjockt på golvetav hennes garderob. De flesta av dem skada fötterna.Få vänner:En kvinna kommer att möta en annan kvinna med gemensamma intressen, göra ett par sakertillsammans, och säga något i stil med "Jag hoppas att vi kan vara goda vänner."En man kommer att möta en annan man med gemensamma intressen, göra ett par sakertillsammans, och säger ingenting. Efter år av att interagera med den här andra mannen,dela förhoppningar och farhågor om att han inte skulle anförtro sig åt sin präst ellerpsykiater, kommer han slutligen svikit sin vakt i ett anfall av berusadsentimentalitet och säga något i stil med "Du vet, för någon som är en sådanryck, jag antar att du är OK. "
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 2desserter:En kvinna i allmänhet beundra ett brokigt dessert för konstnärligarbeta är, prisar sin skapare och väntar en lämplig intervall innanhon motvilligt tar en liten flisa av en kant. En man börjar medta tag i körsbär i centrum.Bil reparation:Den genomsnittliga människan tänker sin Y-kromosom innehåller fullständig reparationmanualer för varje bil som gjorts sedan andra världskriget. Han kommer att arbeta på ett problemsjälv tills det antingen går bort eller förvandlas till något som "inte kan varafast utan specialverktyg ".Den genomsnittliga kvinnan tänker "att roliga dunk-dunk brus" är ennoggrann beskrivning av en bil problem. Hon kommer dock att habil service vid rätt intervall och därmed medföra färre problem änden genomsnittlige mannen.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 4Kläder:Män inte kassera kläder. Den genomsnittliga mannen har fortfarande gymmet skjortanhan bar i high school. Han tror att en jacka är "bara få höggs" omden tid det utvecklar hål i armbågarna. En man kommer att låta nya skjortor sitta påhyllan i sin originalförpackning för ett par år innandem att använda, hoppas de kommer att bli mer bekväm med åldern.Kvinnor tänker kläder är radioaktivt, med en halveringstid på ett år.De utövar försiktighetsåtgärder för att undvika kontaminering av förra årets mode.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 5Förtroende:Den genomsnittliga kvinnan skulle verkligen vilja veta om hennes partner är lurarrunt bakom hennes rygg. Samma kvinna skulle inte berätta för henne bästa vän omhon visste de bästa vänner "mate hade en affär. Hon ska berätta allt henneAndra vänner, dock. Den genomsnittliga mannen kommer inte att säga något om han vet atten av hans väns kompisar lurar runt, och han vill helst inte veta omhans kompis är otrogen heller, av rädsla för att det skulle vara med enav hans vänner. Han kommer att berätta alla sina vänner om sina egna angelägenheter, men,så att de kan vara redo om han behöver ett alibi.Körning:En typisk man tror att han Mario Andretti så snart han glider bakomratten i sin bil. Det faktum att det är en 8-årig Honda håller intehonom från att försöka ut-påskynda killen i Porsche vem försökeratt skära honom; motorväg på ramper är spännande utmaningar att se vem som harRätta virket på morgonen pendla. Har han eller han inte? Endast hans kroppbutik vet säkert. Försäkringsbolagen förstå detta beteende, ochpris sin politik därefter.En kvinna kommer att sakta ner för att låta en bil samman framför henne, och fåbakre slutade med en annan kvinna som var upptagen att lägga sista handen vidhennes makeup.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 6badrum:En man har sex saker i sitt badrum - en tandborste, tandkräm,raklödder, rakhyvel, en bar Dial tvål och en handduk från Holiday Inn.Det genomsnittliga antalet objekt i den typiska kvinnans badrum är 437. En manskulle inte kunna identifiera de flesta av dessa artiklar.Specerier:En kvinna gör en lista över saker som hon behöver och sedan går till affärenoch köper dessa saker. En man väntar 'til de enda objekt kvar i sitt kylskåpär en halv lime och ett blått band. Då han går matinköp. Han köperallt som ser bra ut. Vid tiden som en man når kassadisken,hans vagn packad hårdare att Clampett bil på Beverly Hillbillies.Naturligtvis kommer detta inte att stoppa honom från att komma in i 10-poster eller mindre körfält.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 8Går ut:När en man säger att han är redo att gå ut, betyder det att han är redo att gåut. När en kvinna säger att hon är redo att gå ut, betyder det att hon kommer att vara redoatt gå ut, så snart som hon finner sin örhänge, slutar att sätta på hennes smink,kontroller på barnen, gör ett telefonsamtal till sin bästa vän ...katter:Kvinnor älskar katter. Män säger att de älskar katter, men när kvinnorna inteser, män sparka katter.Avkomma:Ah, barn. En kvinna vet allt om sina barn. Hon vetom tandläkarbesök och fotbollsmatcher och romanser och bästa vänneroch favoritmat och hemliga rädslor och förhoppningar och drömmar. Män är vagtmedveten om några korta människor som bor i huset.
		-- Chamfort

%
FORTUNE Diskuterar Skillnaderna mellan KVINNOR OCH MÄN: # 9Tvätt:Kvinnor tvätta varje par dagar. En man kommer att bära varje artikelkläder han äger, inklusive hans kirurgiska byxor som var hip om åttaår sedan, innan han kommer att göra sitt tvätt. När han är äntligen ur kläder,han kommer att bära en smutsig tröja inifrån och ut, hyra en U-Haul och ta hans bergav kläder till tvättstugan. Män förväntar sig alltid att träffa vackra kvinnor påtvättstugan. Detta är en myt.smeknamn:Om Gloria, Suzanne, Deborah och Michelle träffas för lunch,de kommer att ringa varandra Gloria, Suzanne, Deborah och Michelle. Men omMike, Dave, Rob och Jack gå ut för en Brewsky, de kommer givethänvisa till varandra som Bullet-Head, Godzilla, jordnötter Brain och värdelös.sockor:Män bär förnuftiga strumpor. De bär vanliga vita sweatsocks.Kvinnor bär konstiga strumpor. De skärs långt under anklarna, har bilderav moln på dem, och har en stor luddig boll på baksidan.
		-- Chamfort

%
Fred märkte hans rumskamrat hade en svart öga när han återvände från en dans."Vad hände?""Jag slogs av skönheten i platsen."
		-- Chamfort

%
Vänner var förvånad, faktiskt, när Frank och Jennifer bröt derasengagemang, men Frank hade en klar förklaring: "Vill du gifta sig med någon somvar vanligtvis otrogen, som ljög vid varje tur, som var självisk och latoch sarkastisk? ""Naturligtvis inte", sade en sympatisk vän."Jo", svarade Frank, "varken skulle Jennifer."
		-- Chamfort

%
Från skrivbordet avrapunzelKära Prince:Använd stege i kväll - du dela mina ändar.
		-- Chamfort

%
Äkta lycka är när en kvinna ser en dubbelhaka på sin makesgammal flicka vän.
		-- Chamfort

%
Män är roade av nästan alla idiot sak - det är därför professionella ishockey är så populär - så att köpa presenter till dem är lätt. Men du bordealdrig köpa dem kläder. Män tror att de redan har alla de kläder denågonsin kommer att behöva, och nya gör dem nervösa. Till exempel, din genomsnittligaman har 84 band, men han bär på sin höjd, bara tre av dem. Han har lärt sig,genom förödmjukande försök och misstag, att om han bär någon av de andra 81band, kommer hans fru förmodligen skratta åt honom ( "Du kommer inte att bära denslips med som passar, är du? "). Så han har minskat ner det till tre säkraband, och har gått flera år utan att bli utskrattad. Om du ger honomen ny slips, kommer han att låtsas vilja det, men innerst inne att han kommer att hata dig.Om du vill ge en man något praktiskt, överväga däck. Mer änen gång, skulle jag ha gärna handlas alla gåvor jag fått en ny uppsättning däck.
		-- Dave Barry, "Christmas Shopping: A Survivor's Guide"

%
Flickor snyggare i snöstormar.
		-- Archie Goodwin

%
Flickor gifta för kärlek. Pojkar gifta på grund av en kronisk irritation somfår dem att dras i riktning mot objekt med vissa kroklinjigegenskaper.
		-- Ashley Montagu

%
Flickor egentligen vet precis vad de vill - du räkna ut det själv!
		-- Ashley Montagu

%
Flickor som kastar sig på män, faktiskt tar mycket försiktig mål.
		-- Ashley Montagu

%
Ge en kvinna en tum och hon ska parkera en bil i den.
		-- Ashley Montagu

%
Gud skapade några perfekta huvuden. Resten han täckt med hår.
		-- Ashley Montagu

%
Gud skapade kvinnan. Och tristess har faktiskt upphör från det ögonblicket -men många andra saker upphörde också. Kvinnan var Guds andra misstag.
		-- Nietzsche

%
Bra flickor går till himmel, dåligaflickor går överallt.
		-- Nietzsche

%
Harold hade aldrig ville ha en kvinna så mycket i sitt liv, efter overhearing22-åriga skönheten anmärkning att han var för gammal och ur form för henne. Debestämd septuagenarian inlett omedelbart efter en rigorös självförbättringprogram. Han hade hans ansikte lyft, köpte en tupé, sprang fem miles varje dag,lyfte vikter och antog en strikt vegetarisk kost. Inom några månader, denföryngrad man vann den unga kvinnans hjärta, och hon gick med på att gifta sig med honom.På väg ut ur kapellet, men Harold dödligt slogav blixten. Rasande, konfronterade han Sankte vid pärleporten. "Hurkan du göra så här mot mig efter all smärta jag gick igenom? ""För att vara ärlig, Harold," Saint Peter fåraktigt svarade: "Jag gjorde intekänner igen dig. "
		-- Nietzsche

%
Hatt check flicka:"Godhet Vad vackra diamanter!"Mae West:"Godhet hade ingenting att göra med det, dearie."
		-- "Night After Night", 1932

%
Att ha ett barn är inte så illa. Om du är en kvinnlig kejsare pingvin iAntarktisk. Hon lägger ägg, rullar den över till fadern, sedan tar fartför varmare väder där hon äter och äter och äter. För två månader,far står stel, utan mat, blind i 24-timmars mörk, balanseringägget på fötterna. Efter den lilla pingvinen kläcks, moranser det lämpligt att komma hem.
		-- L. M. Boyd, "Austin American-Statesman"

%
Han gav henne en blick som du kunde ha hälls på en våffla.
		-- L. M. Boyd, "Austin American-Statesman"

%
Den som går in i sin frus omklädningsrum är en filosof eller en dåre.
		-- Balzac

%
Den som är berusad med vin kommer att vara nykter igen i samband mednatt, men han som berusad av munskänken kommer inte återfå sinkänner till dagen för domen.
		-- Saadi

%
Hej, Jim, det är jag, Susie Lillis från tvättstugan. Du sa att du varringer och det har varit två veckor. Vad som är fel, förlorar du mitt nummer?
		-- Saadi

%
Höga klackar är en anordning uppfanns av en kvinna som var trött på att vara kysstepå pannan.
		-- Saadi

%
Honom: "Din hud är så mjuk Är du en modell.?"Hennes: "Nej" [blush] "Jag är en kosmetolog."Honom: "Really Det är otroligt ... Det måste vara mycket svårt att hanteratyngdlöshet. "
		-- "The Jerk"

%
Hans motiv var strikt heder, eftersom uttrycket är: det vill säga, att rånaen dam av hennes förmögenhet i form av äktenskap.
		-- Henry Fielding, "Tom Jones"

%
"Home Sweet Home" måste ju ha skrivits av en ungkarl.
		-- Samuel Butler

%
Horace bästa ode skulle inte tillfredsställa en ung kvinna så mycket som den mediokraverser den unge mannen hon är förälskad i.
		-- Moore

%
Hur mycket för era kvinnor? Jag vill köpa din dotter ... hur mycket förDen lilla tjejen?
		-- Jake Blues, "The Blues Brothers"

%
"Hur skulle jag kunna veta om jag tror på kärlek vid första ögonkastet?" sexigsocial klättrare sade till hennes rumskamrat. "Jag menar, jag har aldrig sett en Porschefull med pengar innan. "
		-- Jake Blues, "The Blues Brothers"

%
Jag är mycket förtjust i sällskap med damer. Jag gillar deras skönhet,Jag gillar deras delikatess, jag gillar deras livlighet, och jag gillar deras tystnad.
		-- Samuel Johnson

%
Jag började för många år sedan, som så många unga män gör, i sökandet efterperfekta kvinnan. Jag trodde att om jag såg tillräckligt länge och hårt nog,Jag skulle hitta henne och då skulle jag vara säker för livet. Tja, åroch romanser kom och gick, och jag så småningom hamnade lösa för någonmycket mindre än min uppfattning om perfektion. Men en dag, efter många årtillsammans, jag låg där på vår säng återhämta sig från en liten sjukdom. Minfru satt på en stol bredvid sängen, surrande mjukt och titta påden sena eftermiddagssolen filtrering genom träden. De enda ljud tillhöras på andra håll var klockan tickar, vattenkokaren nere startatt koka, och en och annan elev passerar under våra fönster. Ochnär jag tittade upp i min fru nu rynkiga ansiktet, men fortfarande varmt ochblinkande ögon, insåg jag något om perfektion ... kommer det baramed tid.
		-- James L. Collymore, "Perfect Woman"

%
Jag tror att en liten inkompatibilitet är livets krydda, särskilt om hanhar inkomster och hon är pattable.
		-- Ogden Nash

%
Jag kan känna för henne eftersom, även om jag aldrig har varit en Alaskan prostitueraddansar på baren i en spangled klänning, jag fortfarande får mycket uttråkad med tvättoch strykning och disk och matlagning dag efter obevekliga dag.
		-- Betty MacDonald

%
Jag kan inte para sig i fångenskap.
		-- Gloria Steinem, on why she has never married.

%
Jag kommer från en liten stad vars befolkning aldrig ändrats. Varje gång en kvinnablev gravid, någon lämnat staden.
		-- Michael Prichard

%
Jag njuta av en god lång promenad - särskilt när min fru tar en.
		-- Michael Prichard

%
"Jag behöver inte ta detta missbruk från dig - jag har hundratalsmänniskor väntar på att missbruka mig. "
		-- Bill Murray, "Ghostbusters"

%
Jag antar att jag aldrig glömma henne. Och kanske jag inte vill. hennes andevar vild, som en vild apa. Hennes skönhet var som en vacker hästrids av en vild apa. Jag glömmer hennes andra kvaliteter.
		-- Jack Handey, The New Mexican, 1988.

%
Jag har svårt att bli attraherad av någon som kan slå mig.
		-- John McGrath, Atlanta sportswriter, on women weightlifters.

%
Jag har funnit det omöjligt att bära den tunga bördan av ansvar ochatt fullgöra mina plikter som kung som jag skulle vilja göra utan hjälp ochstöd för kvinnan jag älskar.av den brittiska tronen för att gifta sig med den amerikanskafrånskild Wallis Warfield Simpson.
		-- Edward, Duke of Windsor, 1936, announcing his abdication

%
Jag har nu kommit fram till att aldrig mer tänka på att gifta sig,och av denna anledning: Jag kan aldrig vara nöjd med någon som skullevara dumskalle nog att ha mig.
		-- Abraham Lincoln

%
Jag vet placeringen av kvinnor: när du kommer, kommer de inte; närdu kommer inte, sätter de sina hjärtan på er egen lutning.
		-- Publius Terentius Afer (Terence)

%
Jag lärde mig att spela gitarr bara för att få flickor och alla som säger att deinte bara ljuger!
		-- Willie Nelson

%
Jag gillar att vara singel. Jag är alltid där när jag behöver mig.
		-- Art Leo

%
Jag gillar mig, men jag kommer inte att säga att jag är så vacker som tjuren som kidnappadeEuropa.
		-- Marcus Tullius Cicero

%
Jag gillar unga flickor. Deras berättelser är kortare.
		-- Tom McGuane

%
Jag älskar att vara gift. Det är så stor att finna att en speciell persondu vill irritera för resten av ditt liv.
		-- Rita Rudner

%
Jag älskar Mickey Mouse mer än någon kvinna jag någonsin känt.
		-- Walt Disney

%
Jag lyckades att säga "Sorry" och inget mer. Jag visste att han ogillademig att gråta.Den här gången sade han tittar på mig, "Vid vissa tillfällen är det bättreatt gråta."Jag lägger mitt huvud på bordet och snyftade: "Om bara hon kunde kommatillbaka; Jag skulle vara trevligt. "Francis sade: "Du gav henne stort nöje alltid.""Åh, inte tillräckligt.""Ingen kan ge någon tillräckligt."	"Aldrig?""Nej, inte alltid. Men man måste gå på att försöka.""Och inte någonsin värderar människor tills de är borta?""Sällan", sade Francis. Jag gick på gråt; Jag såg hur lite jag hadevärderas honom; hur lite jag hade värderat något som var mitt.
		-- Pamela Frankau, "The Duchess and the Smugs"

%
Jag gifte under mig. Alla kvinnor gör.
		-- Lady Nancy Astor

%
Jag träffade en underbar ny människa. Han är fiktiv, men du kan inte få allt.
		-- Cecelia, "The Purple Rose of Cairo"

%
Jag har aldrig förväntas se den dag då flickor skulle få solbrända iplatser de gör idag.
		-- Will Rogers

%
Jag har aldrig träffat en kvinna som jag inte kunde dricka söt.
		-- Will Rogers

%
Jag läste Playboy av samma anledning jag läste National Geographic. Att sesevärdheterna Jag kommer aldrig att besöka.
		-- Will Rogers

%
Jag vägrar att förpassa hela manligt kön till plantskolan. Jag insisterar påtro att vissa män är mina jämlikar.
		-- Brigid Brophy

%
Jag respekterar äktenskapet som institution. Jag har alltid trott att varjekvinna ska gifta sig - och ingen människa.
		-- Benjamin Disraeli, "Lothair"

%
Jag satt bredvid henne, sa hej, erbjöd sig att köpa henne en drink ... och sedannaturligt urval uppfödda sitt fula huvud.
		-- Benjamin Disraeli, "Lothair"

%
Jag tror att hon måste ha varit mycket strikt uppfostrad, hon är så desperatangelägna om att göra fel sak på rätt sätt.
		-- Saki, "Reginald on Worries"

%
Jag tror att världen är redo för historien om en ful ankunge som växte upp tillförbli en ful ankunge, och levde lyckliga i alla sina dagar.
		-- Chick

%
Jag vill köpa en make som varje vecka när jag sitter ner för att titta "St.På andra håll ", inte kommer att skrika," Glöm det, Blanche ... Det är dags för Hee-Haw! "
		-- Berke Breathed, "Bloom County"

%
Jag vill gifta sig med en flicka precis som flickan som gift kära gamla pappa.
		-- Freud

%
Jag var i en skönhetstävling en. Jag inte bara kom i förra var jag slog imunnen av Miss Secret Agent.
		-- Phyllis Diller

%
Jag var inte kyssa henne, jag viskade i hennes mun.
		-- Chico Marx

%
Jag kommer inte att säga att kvinnor har inget tecken; snarare, de har en nyen varje dag.
		-- Heine

%
Jag skulle gärna höja min röst i beröm av kvinnor, bara de inte kommer att låta mighöja min röst.
		-- Winkle

%
Jag skulle inte gifta sig med henne med en tio fot stolpe.
		-- Winkle

%
Jag skulle nog nöja sig med en vampyr om han var tillräckligt romantisk.Det gick inte att vara något sämre än några av de relationer som jag har haft.
		-- Brenda Starr

%
Jag vill hellre ha två flickor vid 21 var än en flicka på 42.
		-- W. C. Fields

%
Jag försvarar hennes ära, vilket är mer än hon någonsin gjort.
		-- W. C. Fields

%
Jag är inte denyin "kvinnorna är dåraktig: Gud Allsmäktig gjort dem att matcha män.
		-- George Eliot

%
Jag är väldigt gammaldags. Jag tror att människor ska gifta sig för livet,som duvor och katoliker.
		-- Woody Allen

%
Jag har varit i flera varv än en servett.
		-- Mae West

%
Jag har tillbringat nästan hela mitt liv med mycket intelligenta män. Dom är inteliksom andra män. Deras ande är stor och stimulerande. De hatar strid;ja de avvisar det. Deras uppfinningsrika gåvor är gränslös. de kräverhängivenhet och lydnad. Och en känsla för humor. Jag lyckligtvis gav allt detta.Jag hade tur att väljas och smart nog att förstå dem.
		-- Marlene Dietrich, on her friendship with Ernest Hemingway

%
Om jag var tvungen att leva mitt liv igen, skulle jag göra samma misstag, bara förr.
		-- Tallulah Bankhead

%
Om jag sa att du hade en vacker kropp, skulle du håller den mot mig?
		-- Tallulah Bankhead

%
Om det inte vore för de presenter, skulle en rymning vara att föredra.
		-- George Ade, "Forty Modern Fables"

%
Om män agerade efter äktenskapet som de gör under uppvaktning, det skullefärre skilsmässor - och fler konkurser.
		-- Frances Rodman

%
Om någon skulle fråga mig för en genväg till sensualitet, skulle jagföreslår han gå och handla för en begagnad 427 Shelby-Cobra. Men det är bararättvist att varna dig om att av de 300 män som bytte till dem 1966,bara två gick tillbaka till kvinnor.
		-- Mort Sahl

%
Om flickan du älskar flyttar in med en annan kille en gång, det är mer än tillräckligt.Två gånger, det är alldeles för mycket. Tre gånger, det är historien om ditt liv.
		-- Mort Sahl

%
Om det finns någon realistisk avskräckande för äktenskap, är det faktum att duhar inte råd skilsmässa.
		-- Jack Nicholson

%
Om vi ​​män gifte de kvinnor vi förtjänade, skulle vi ha en mycket dålig tid för det.
		-- Oscar Wilde

%
Om kvinnor ska vara mindre rationella och mer emotionella påi början av vår menstruationscykeln, när det kvinnliga könshormonet är somlägsta nivå, varför är det inte logiskt att säga att i dessa få dagarkvinnor beter mest som hur män beter hela månaden?
		-- Gloria Steinham

%
Om kvinnor inte existerade, skulle alla pengar i världen har ingen betydelse.
		-- Aristotle Onassis

%
Om du är rädd för ensamheten, inte gifta sig.
		-- Anton Chekhov

%
Om du letar efter ett vänligt, well-to-do äldre herre som är ingenlängre intresserad av sex, ta ut en annons i The Wall Street Journal.
		-- Abigail Van Buren

%
Om du ger en man nog rep, kommer han hävdar att han är bunden på kontoret.
		-- Abigail Van Buren

%
Om du gifta sig med en man som är otrogen mot sin fru, kommer du vara gift med en man somotrogen mot sin fru.
		-- Ann Landers

%
Om du måste gifta, är det alltid klokt att gifta sig med skönhet.Annars kommer du aldrig att hitta någon att ta bort henne händerna.
		-- Ann Landers

%
Om du vill att jag ska vara en bra liten kanin bara dingla några karat framförnäsan.
		-- Lauren Bacall

%
Om du vill bli förstört, gifta sig med en rik kvinna.
		-- Michelet

%
Om du vill läsa om kärlek och äktenskap du har att köpa två separataböcker.
		-- Alan King

%
Om du vill att din make att lyssna och betala strikt uppmärksamhet åt varjeord du säger, tala i sömnen.
		-- Alan King

%
Om du vill kvinnor att älska dig, vara original; Jag känner en man som bar pälsstövlar sommar och vinter, och kvinnorna blev kär i honom.
		-- Anton Chekhov

%
Att köpa hästar och ta en hustru blunda tätt och lovordarsjälv till Gud.
		-- Anton Chekhov

%
I kristendomen kan en man ha endast en hustru. Detta kallas monotoni.
		-- Anton Chekhov

%
I äktenskap, som i krig, är det tillåtet att ta varje fördel av fienden.
		-- Anton Chekhov

%
I äldre tider offer gjordes vid altaret - en praxis som ärfortfarande fortsatte.
		-- Helen Rowland

%
Mitt i en av de vildaste parterna han någonsin hade varit till den unge mannenmärkt en mycket prydligt och vacker flicka sitta tyst bortsett från resten avfestprissar. Närmar henne, presenterade han sig och efter en tystkonversation, sade: "Jag är rädd att du och jag inte riktigt passar in i dettaavtrubbad grupp. Varför jag inte ta dig hem? """Fine", sa flickan, leende upp på honom demurely. "Var bor du?"
		-- Helen Rowland

%
Insanity anses vara en grund för skilsmässa, men av sammatoken är det kortaste avstickare till äktenskap.
		-- Wilson Mizner

%
Är ett bröllop lyckas om det lossnar utan problem?
		-- Wilson Mizner

%
Är inte äktenskapet en öppen fråga, när det påstås, frånbörjan av världen, att sådana som är i institutet vill fåut, och som är ute vill komma in?
		-- Ralph Emerson

%
Är det inte ironiskt att många män tillbringar en stor del av deras livundvika äktenskap medan målmedvetet driva de saker somskulle göra dem bättre framtidsutsikter?
		-- Ralph Emerson

%
Det [äktenskapet] händer som med burar: fåglarna utan förtvivlanatt komma in, och de inom förtvivlan av att få ut.
		-- Michel Eyquem de Montaigne

%
Det förekom inte att min varelse med två män kontinuerligt skulleränta någon eller väcka någons betänkligheter. Jag bad om en inbjudanför Heinrich också, så ofta som det verkade möjligt, när Paulus och jag varinbjuden till ett samkväm. Jag kände uppsättning regler andra levde medvar irrelevant. Min barndom inställning - varje försök att justera ärhopplös och du kan lika gärna följa dina egna attityder - måste habar mig.
		-- Hannah Tillich, "From Time to Time"

%
Det är inte mycket beteckna som ett gifter, för en är säker på att hitta utNästa morgon var det någon annan.
		-- Will Rogers

%
Det har med rätta observerats av vise i alla länder att även om en människa kan varamest lyckligt gift och fortsätter i detta tillstånd med största belåtenhet,det inte nödvändigtvis att han har därför slagit stenblinda.
		-- H. Warner Munn

%
Det är alltid bättre att besöka hem med en vän. Dina föräldrar kommerinte vara nöjd med denna plan, eftersom de vill att ni alla för sig själva ocheftersom det i närvaro av en vän, måste de agera som mognamänniskor.Den värsta sortens vän att ta hem är en flicka, för i så fall,det finns potential att dina föräldrar kommer att förlora dig inte bara förvaraktighet besök men alltid. Den värsta sortens flicka att ta hem är enav en annan religion: Inte bara kommer du att gå förlorade till dina föräldrar alltid mendu kommer att gå förlorade till en kvinna som är immun mot deras religiösa / moraliska argumentoch vars exempel kommer oåterkalleligen korrupta dig.Låt oss säga att du har blivit kär i just en sådan flicka och villatt ta henne hem för semester. Du är medveten om dina föräldrars främlingsfientligsvar på någon av en annan religion. Hur man förbereder dem för chocken?Enkelt. Kalla dem strax innan ditt besök och berätta att duhar blivit ganska allvarligt om någon som är av en annan religion, enannan ras och samma kön. Säg att du redan har anmodatperson att möta dem. Ge informationen en stund att sjunka in och sedanpåpeka att du bara skojade, att din älskare är bara en annanreligion. De kommer att bli så lättad att de kommer att välkomna henne med öppna armar.
		-- Playboy, January, 1983

%
Det förklaras att alla relationer kräver lite givande och tagande. Dettaär osant. Alla partnerskap kräver att vi ger och ger och ger och påsist, när vi floppar i våra gravar utmattad, får vi veta att vi inte gavtillräckligt.
		-- Quentin Crisp, "How to Become a Virgin"

%
Det är meningslöst att försöka prata en ung kvinna ur hennes passion:kärlek ligger inte i örat.
		-- Walpole

%
Det är de farligaste idag för en man att betala någon uppmärksamhet till hansfru offentligt. Det gör alltid människor tror att han slår henne närde är ensamma. Världen har blivit så misstänksam mot något som sersom ett lyckligt gift liv.
		-- Oscar Wilde

%
Det är inte nödvändigt att undersöka huruvida en kvinna vill ha något fördessert. Svaret är ja, hon vill ha något för dessert, menHon skulle vilja att ni beställa det så att hon kan ta på det med din gaffel. Honinte vill att du ska uppmärksamma detta genom att säga: "Om du ville ha endessert, varför inte du beställer en? " Du måste förstå, hon hardessert hon vill. Dessert hon vill är innesluten i din.
		-- Merrill Markoe, "An Insider's Guide to the American Woman"

%
Det är nu helt lagligt för en katolsk kvinna att undvika graviditet genom en utväg attmatematik, även om hon fortfarande förbjudet att ta till fysik och kemi.
		-- H. L. Mencken

%
Det är möjligt att blondiner föredrar också herrar.
		-- Maimie Van Doren

%
Det tar en smart man att ha sista ordet och inte använda den.
		-- Maimie Van Doren

%
Det var en fin, söt natt, den trevligaste sedan min skilsmässa, kanske finastesedan mitten av mitt äktenskap. Det fanns energi, mjukhet, nåd ochskratt. Jag tog även mina strumpor. I min cirkel, betyder den klassen.
		-- Andrew Bergman "The Big Kiss-off of 1944"

%
Det regnade kraftigt, och bilisten hade problem med bilen på en ensam landväg. Angelägna om att hitta tak över huvudet för natten, gick han över till en bondgårdoch knackade på ytterdörren. Ingen svarade. Han kunde känna vattnetfrån taket löper längs nacken när han stod på farstubron.Nästa gång han knackade högre, men fortfarande inget svar. Vid det här laget var han indränkttill huden. Desperat han krossas på dörren. Äntligen huvudet av enman dök upp i en övervåningen fönster.	"Vad vill du?" frågade han buttert."Min bil gick sönder", sade resenären, "och jag vill veta om duskulle låta mig stanna här för natten. ""Visst", svarade mannen. "Om du vill stanna kvar hela natten, är detokej med mig. "
		-- Andrew Bergman "The Big Kiss-off of 1944"

%
Det var inte precis en skilsmässa - Jag handlades.
		-- Tim Conway

%
Det är en rolig sak som när en kvinna inte har fått någotpå jorden för att oroa sig för, går hon bort och gifter sig.
		-- Tim Conway

%
"Det är män som han som ger Y-kromosomen ett dåligt rykte."
		-- Tim Conway

%
Det är inte initialt kjol längd, det är upcreep.
		-- Tim Conway

%
Det är inte män i mitt liv, men livet i mina män som räknas.
		-- Mae West

%
Det är bra tjejer som håller dagböcker, dåliga flickor aldrig har tid.
		-- Tallulah Bankhead

%
Det är teorin om Jess Birnbaum, av Time magazine, att kvinnor meddåliga ben bör hålla sig till långa kjolar, eftersom de täcker en mängd smalbenen.
		-- Tallulah Bankhead

%
Joe satt som sin döende hustrus säng.Hennes röst var lite mer än en viskning."Joe, älskling", säger hon andades, "Jag har en bekännelse att görainnan jag går. Jag ... Jag är en som tog $ 10.000 från din säkra ...Jag tillbringade det på en fling med din bästa vän, Charles. Och det var jag somtvingade din älskarinna att lämna staden. Och jag är den som rapporteradedin inkomst skatteflykt till I.R.S ... ""Det är okej, kära, inte ge det en andra tanke,"viskade Joe. "Jag är en som förgiftade dig."
		-- Tallulah Bankhead

%
Precis som jag inte kan minnas någon tid när jag inte kunde läsa och skriva, jag kan inteminns helst när jag inte utöva min fantasi i dagdrömmar omkvinnor.
		-- George Bernard Shaw

%
Kath: Kan han vara närvarande vid födseln av sitt barn?Ed: Det är någon rimlig barn kan förvänta sig om pappa är närvarandevid befruktningen.
		-- Joe Orton, "Entertaining Mr. Sloane"

%
Föra dagbok och en dag kommer att hålla dig.
		-- Mae West

%
Håll kvinnor du inte kan. Gifta sig med dem och de kommer att hata hur du gårtvärs över rummet; förblir deras älskare, och de jilt dig i slutet av sexmånader.
		-- Moore

%
Håll ögonen vidöppna före äktenskapet, halv stänga efteråt.
		-- Benjamin Franklin

%
Kyssa din hand kan göra dig mycket bra, men en diamant ochsafir armband varar för evigt.
		-- Anita Loos, "Gentlemen Prefer Blondes"

%
Lady Nancy Astor:"Winston, om du var min man, jag skulle sätta gift i ditt kaffe."Winston Churchill:"Nancy, om du var min fru, jag skulle dricka det."
		-- Anita Loos, "Gentlemen Prefer Blondes"

%
Lank: Här går vi. Vi håller på att sätta ett nytt rekord.Earl: (till publiken) Vad sägs om ett datum?Lank: Vi har gjort det. Earl har satt ett nytt rekord. Avvisades av      20.000 kvinnor.
		-- Lank and Earl

%
Stora ökningar i kostnader med tvivelaktiga ökningar i prestanda burktolereras endast i kapplöpningshästar och kvinnor.
		-- Lord Kelvin

%
Låt din piga tjänare vara trogen, stark och hemtrevlig.
		-- Benjamin Franklin

%
Låt oss bara säga att när en förändring krävdes, justerade jag. i varjerelation som existerar, människor måste söka ett sätt att överleva. om duverkligen bryr sig om personen du göra vad som krävs, eller är det slut.För första gången, fann jag att jag verkligen skulle kunna ändra och egenskaperJag mest beundrade i mig själv jag gav upp. Jag slutade vara högt och diktatorisk ...Åh, okej. Jag var fortfarande högt och diktatorisk, men bara bakom ryggen.
		-- Kate Hepburn, on Tracy and Hepburn

%
Livet börjar vid mittuppslag och expanderar utåt.
		-- Miss November, 1966

%
Livet i det här samhället är, i bästa fall, en fullkomlig hål och ingen aspekt av samhälletatt alls relevant för kvinnor, det återstår att medborgerligt sinnade ansvarigspänningssökande kvinnor endast att störta regeringen, eliminera pengarsystemet, institut fullständig automatisering och förstöra det manliga könet.
		-- Valerie Solanas

%
Livet suger. Cynisk, människofientliga manlig, 34, letar efter själsfrände, menvissa inte att hitta henne. Släpp mig en anteckning. Jag ringer dig, kommer vi att tala ochJag kommer att be dig på middag där jag kommer förmodligen tillbringar mer än jag kanråd i ett svagt försök att imponera på dig. Sedan kommer vi att inse att vi harabsolut ingenting gemensamt och vi kommer att gå skilda vägar, merförbittrade och deprimerad än tidigare (om något sådant är möjligt).
		-- Valerie Solanas

%
Livet är för kort för att dansa med fula kvinnor.
		-- Valerie Solanas

%
Liksom alla unga män, du kraftigt överdriver skillnaden mellan enung kvinna och en annan.
		-- George Bernard Shaw, "Major Barbara"

%
Liksom skidorten flickor söker män och män som sökerför flickor, är situationen inte så symmetrisk som det kan tyckas.
		-- Alan McKay

%
Små flickor, som fjärilar, behöver ingen ursäkt.
		-- Lazarus Long

%
Ensamma män söker sällskap. Ensamma kvinnor sitta hemma och vänta.De träffas aldrig.
		-- Lazarus Long

%
Massor av flickor kan fås för en låt. Tyvärr, ofta visar det sig attär det bröllopsdagen marsch.
		-- Lazarus Long

%
Kärlek är en idealisk sak, äktenskapet en real thing; en sammanblandning av den verkligamed den ideala aldrig går ostraffade.
		-- Goethe

%
Kärlek är en tvångsmässig illusion som botas genom äktenskap.
		-- Dr. Karl Bowman

%
Kärlek är villfarelsen att en kvinna skiljer sig från en annan.
		-- H. L. Mencken

%
Kärleken gör dumbommar, äktenskap cuckolds och patriotism illvilliga idioter.
		-- Paul Leautaud, "Passe-temps"

%
Macho bevisar inte mucho.
		-- Zsa Zsa Gabor

%
Man och hustru gör en dåre.
		-- Zsa Zsa Gabor

%
Mången har blivit kär i en flicka i en ljus så mörk att han skulleinte ha valt en kostym av den.
		-- Maurice Chevalier

%
Mången kär i en grop gör misstaget att gifta sigHela flicka.
		-- Stephen Leacock

%
Många en man som tror att han kommer på en jungfrufärd meden kvinna får reda på senare att det var bara en shake-down kryssning.
		-- Stephen Leacock

%
Många fru tror att hennes make är världens största älskare.Men hon kan aldrig fånga honom på det.
		-- Stephen Leacock

%
Många män gå sönder på pengarna deras fruar spara på försäljningen.
		-- Stephen Leacock

%
Äktenskap alltid kräver den största förståelse för konsten attinsincerity möjligt mellan två människor.
		-- Vicki Baum

%
Äktenskap orsakar dejting problem.
		-- Vicki Baum

%
Äktenskapet är en hemsk offentlig bekännelse av en strikt privat avsikt.
		-- Vicki Baum

%
Äktenskapet är en stor institution - men jag är inte redo för en institution ännu.
		-- Mae West

%
Äktenskapet är en mycket som armén, klagar alla, men du skulle varaförvånad över det stora antal som åter värva.
		-- James Garner

%
Äktenskapet är en roman där hjälten dör i det första kapitlet.
		-- James Garner

%
Äktenskapet är en tre ring cirkus: förlovningsring, vigselring, och lidande.
		-- Roger Price

%
Äktenskapet är en institution där två åtar sig att bli en och enförbinder sig att bli någonting.
		-- Roger Price

%
Förbindelse är baserad på teorin att när en man upptäcker ett märke av ölexakt hans smak han skulle genast kasta upp sitt jobb och gå till jobbeti bryggeriet.
		-- George Jean Nathan

%
Äktenskapet är att lära sig om kvinnor den hårda vägen.
		-- George Jean Nathan

%
Äktenskapet är som snurrar en stafettpinne, vrida handsprings eller äta medpinnar. Det ser lätt tills du prova det.
		-- George Jean Nathan

%
Äktenskapet är lågt, men du tillbringa resten av ditt liv att betala för det.
		-- Baskins

%
Äktenskapet är inte bara dela fettucine, men delabördan av att finna fettucine restaurangen i första hand.
		-- Calvin Trillin

%
Förbindelse är den enda äventyr öppna för feg.
		-- Voltaire

%
Äktenskapet är en process för att ta reda på vilken typ av människa din fru skulleha föredragit.
		-- Voltaire

%
Äktenskapet är papperskorgen av känslor.
		-- Voltaire

%
Äktenskap, i livet, är som en duell mitt i en strid.
		-- Edmond About

%
Äktenskap görs i himlen och fullbordade på jorden.
		-- John Lyly

%
Gifta sig i hast och alla börjar räkna månaderna.
		-- John Lyly

%
Äktenskapet är roten till allt ont.
		-- John Lyly

%
Äktenskapet är inte ett ord, det är en mening.
		-- John Lyly

%
Män är alltid redo att respektera något som tråkar ut dem.
		-- Marilyn Monroe

%
Män är de varelser med två ben och åtta händer.
		-- Jayne Mansfield

%
Män är inte attraherad av mig genom mitt sinne. De lockas av vad jaginte har något emot ...
		-- Gypsy Rose Lee

%
Män har en mycket bättre tid det än kvinnor; för en sak de gifter sig senare;för en annan sak som de dör tidigare.
		-- H. L. Mencken

%
Män har som överdrivna en uppfattning om sina rättigheter som kvinnor har sina fel.
		-- E. W. Howe

%
Män lever för tre saker, snabba bilar, snabba kvinnor och snabbmat.
		-- E. W. Howe

%
Män gör aldrig passerar på flickor som bär glasögon.
		-- Dorothy Parker

%
Män kvalitet är inte rädda för kvinnor för jämställdhet.
		-- Dorothy Parker

%
Män säger kvinnor vad behagar dem; kvinnor gör med män vad som behagar dem.
		-- DeSegur

%
Män visar sällan gropar till flickor som har finnar.
		-- DeSegur

%
Män minns fortfarande den första kyssen efter kvinnor har glömt den sista.
		-- DeSegur

%
Män som omhuldar för kvinnor högsta respekt är sällan populärt med dem.
		-- Joseph Addison

%
Herrtidningar har ofta bilder på nakna damer. Damtidningarockså ofta har bilder på nakna kvinnor. Detta beror på att den kvinnligakropp är en vacker konstverk, medan den manliga kroppen är hårig och knottrig ochbör inte ses av dagens ljus.
		-- Richard Roeper, "Men and Women Are Different"

%
Miguel Cervantes skrev Donkey Hote. Milton skrev Paradise Lost, då hanshustru dog och han skrev Paradise återfått.
		-- Richard Roeper, "Men and Women Are Different"

%
Moe: Wanna spela poker i kväll?Joe: Jag kan inte. Det är barnens utekväll.Moe: Så?Joe: Jag måste stanna hemma med sjuksköterskan.
		-- Richard Roeper, "Men and Women Are Different"

%
Moe: Vad gav du din fru för Alla hjärtans dag?Joe: Den vanliga gåva - hon åt mitt hjärta.
		-- Richard Roeper, "Men and Women Are Different"

%
Pengar och kvinnor är de mest eftertraktade och minst kända av tvåsaker som vi har.
		-- The Best of Will Rogers

%
Pengar är en kraftfull afrodisiakum. Men blommor fungerar nästan lika bra.
		-- Lazarus Long

%
Monogami är den västerländska sed en fru och knappt några älskarinnor.
		-- H. H. Munro

%
... De flesta av oss lärt sig om kärlek den hårda vägen. Även varningar är förmodligenvärdelös, för på något sätt, trots de svåraste varningar om föräldrar och vänner,hundratals har tusentals kvinnor glömt sig i sista minutenoch dukade under för lögner, löften, smicker, eller bara uppmärksamhet avlusting, vackra män, landar sig i komplicerade predikament frånsom en del av dem aldrig återhämtat sig under hela sitt liv. Och jag är intetalar bara dina tonårs Midwesterners 1958; Jag talar om kvinnorav alla åldrar i varje stad i varje år. Den ökända sexuella revolutionenhar räddat ingen från smärta och förvirring av kärlek.
		-- Alix Kates Shulman

%
Min uppfattning om en man vid fyrtio är att en kvinna ska kunna ändra honom,som en sedel, för två tjugoårsåldern.
		-- Alix Kates Shulman

%
Aldrig acceptera en inbjudan från en främling om han ger dig godis.
		-- Linda Festa

%
Aldrig argumentera med en kvinna när hon är trött - eller vilade.
		-- Linda Festa

%
Aldrig äta på en plats som heter mammas. Spela aldrig kort med en man vid namn Dok.Och aldrig ligga ner med en kvinna som har fått mer bekymmer än du.
		-- Nelson Algren, "What Every Young Man Should Know"

%
Aldrig gå till sängs arg. Stanna upp och slåss.
		-- Phyllis Diller, "Phyllis Diller's Housekeeping Hints"

%
Aldrig sova med en kvinna vars problem är värre än din egen.
		-- Nelson Algren

%
berättar aldrig. Inte om du älskar din fru ... Faktum är att om din gamla dam promenaderin på dig, förneka det. Ja. Bara platta ut och hon ska tro det: "Jag ärTellin 'ya. Den här tjejen kom ner med en skylt runt halsen `LayOvanpå mig eller ska jag dör ". Jag visste inte vad jag skulle göra ... "
		-- Lenny Bruce

%
Nyårsafton är den tid på året då en man mest känner hans ålder,och hans hustru påminner oftast honom att handla det.
		-- Webster's Unafraid Dictionary

%
Ingen vänskap är så hjärtlig eller så läcker som för flicka för flicka;inget hat så intensiv eller fast som för kvinnan för kvinnan.
		-- Landor

%
Ingen människa kan ha en rimlig uppfattning av kvinnor tills han länge har förloratintresse hårväxt.
		-- Austin O'Malley

%
Ingen modern kvinna med en nypa känsla någonsin skickar små lappar till enogift man - inte förrän hon är gift, i alla fall.
		-- Arthur Binstead

%
Ingen vet som en kvinna hur man säger saker som är på gång mild och djup.
		-- Hugo

%
Ingen self-made man någonsin gjorde ett så bra jobb som någon kvinna intevill göra några ändringar.
		-- Kim Hubbard

%
Ingen kvinna kan kalla sig fri tills hon kan välja medvetet omhon kommer eller inte kommer att vara en mor.
		-- Margaret H. Sanger

%
Ingen kvinna kan uthärda ett spel man, om han är en stadig vinnare.
		-- Lord Thomas Dewar

%
Ingen kvinna någonsin blir kär i en man om hon har en bättre uppfattning avhonom än han förtjänar.
		-- Edgar Watson Howe

%
Ingen vet riktigt vad lycka är, tills de är gifta.Och då är det för sent.
		-- Edgar Watson Howe

%
Inte alla problem någon har med sin flickvän är nödvändigtvis beror pådet kapitalistiska produktionssättet.
		-- Herbert Marcuse

%
Av alla djur, är pojken mest ohanterliga.
		-- Plato

%
Naturligtvis en platonisk relation är möjligt - men endast mellanman och hustru.
		-- Plato

%
När en kvinna har givit dig hennes hjärta kan man aldrig bli av med resten av henne.
		-- Vanbrugh

%
En gång i tiden fanns det en vacker ung flicka med en promenadgenom skogen. Allt på en gång hon såg en extremt ful tjur groda sittandepå en stock och hennes förvåning grodan talade till henne. "Maiden" kraxade dengroda, "skulle du göra mig en tjänst? Det kommer att bli svårt för dig att tro, menJag var en gång en vacker, charmig prins och sedan ett medelvärde, fula gamla häxan casten stava över mig och vände mig till en groda. ""Åh, vad synd!", Utbrast flickan. "Jag ska göra allt jag kan för atthjälper dig att bryta en sådan spell. ""Jo", svarade grodan "det enda sättet att denna formel kan varatas bort är för vissa vacker ung kvinna att ta mig hem och låt mig spenderanatten under kudden. "Den unga flickan tog fula groda hem och placerade honom under hennekudde på natten när hon gick i pension. När hon vaknade nästa morgon, säkernog finns bredvid henne i sängen var en mycket ung, stilig man, uppenbarligen avkungligt blod. Och så levde de lyckliga i alla sina dagar, förutom att denna daghennes far och mor fortfarande inte tror hennes berättelse.
		-- Vanbrugh

%
En gång i tiden fanns det tre bröder som var riddarepå ett visst rike. Och, det fanns en Princess i ett angränsande rikesom var i giftasvuxen ålder. Tja, en dag, i full rustning, deras hästar,och deras sida, de tre bröderna iväg för att se om någon av dem kundevinna handen. Vägen var lång och det fanns många hinder påsätt, rånare som måste övervinnas, hård terräng att passera. När de klaratvarje hinder de blev mer och mer äcklad av deras sida. Han varinte bara oduglig, var han feg, kunde han inte hantera hästarna, var han,kort sagt, en komplett flopp. När de anlände till domstolen i riket,De fann att de förväntas presentera prinsessan med någraskatt. De två äldre bröder avskräckt, eftersom de inte hadetänkt på detta och var oförberedd. Den yngsta, men hadesvara: Lova henne något, men ge henne vår sida.
		-- Vanbrugh

%
En kväll talade han. Sitter vid hennes fötter, hans ansikte höjas till henne,han lät sin själ att höras. "Min älskling, vad du vill, vad som helstJag är allt jag någonsin kan vara ... Det är vad jag vill erbjuda dig - intesaker som jag får för dig, men saken i mig som gör mig kunna fådem. Det där - man kan inte avstå från det - men jag vill avstå från det - såatt det kommer att bli din - så att det kommer att vara i din tjänst -. endast för dig "Flickan log och frågade: "Tror du jag är sötare än MaggieKelly? "Han fick upp. Han sade ingenting och gick ut ur huset. han aldrigsåg att flickan igen. Gail Wynand, som berömde sig på aldrig behöver enlektion två gånger, inte bli kär igen i åren som följde.
		-- Ayn Rand, "The Fountainhead"

%
En flicka kan vara ganska - men ett dussin är bara en kör.
		-- F. Scott Fitzgerald, "The Last Tycoon"

%
Man föds inte en kvinna, man blir en.
		-- Simone de Beauvoir

%
En mans dårskap är en annan mans hustru.
		-- Helen Rowland

%
Man bör alltid vara kär. Det är anledningen bör man aldrig gifta sig.
		-- Oscar Wilde

%
Endast två grupper av människor faller för smicker - män och kvinnor.
		-- Oscar Wilde

%
Människor i alla typer av kön rapporterar stora svårigheter,dessa dagar, att välja rätt ord att hänvisa till dem av den kvinnligaövertalning."Lady", "kvinna" och "flicka" är alla helt bra ord, menfelaktig tillämpning dem kan tjäna en något från ansvar för vulgaritet till en braswift smack. Vi Messing här med frågor om respekt, nedlåtenhet,respekt, bigotteri, och två vaga begrepp, ålder och rang. Det är oroandetillräckligt för att få raka som är verkligen vad. De som medvetet missbrukarvillkoren i en misbegotten försök till smicker ber om det.En kvinna är någon vuxen kvinnlig person. En flicka är FN-vuxenversion. Om du ringer en pissa sak med knubbiga kinder och rosa hårband en"Kvinna" kommer du förmodligen inte hamnar i trubbel, och om du gör, kommer du attkunna hantera det eftersom hon kommer att vara under tre fot lång. Men om dukallar en vuxen med ett barns namn för den skull innebär att hon har enungdomlig kropp, är du också innebär att hon har en hjärna för att matcha.
		-- Oscar Wilde

%
Fysiskt finns det ingenting att skilja det mänskliga samhället frångård gård förutom att barn är mer besvärligt och kostsamt änkycklingar och kvinnor är inte så helt förslavade som gården lager.
		-- George Bernard Shaw, "Getting Married"

%
Rika ungkarlar bör beskattade. Det är inte rättvist att vissa mänbör vara lyckligare än andra.
		-- Oscar Wilde

%
Sally: C'mon, Ted, allt jag ber dig att göra är att dela dina känslor	med mig.Ted: ALL? Inser du vad du frågar? Män är inte utbildade	att dela. Vi är utbildade för att skydda oss själva genom att intelåta någon för nära. Bra sorg, om jag går runtdela allt med dig, kan du hänga mig på tork.Sally: Den heter "förtroende", Ted.Ted: "Dela"? "Förtroende"? Du verkligen ber mig att segla inokända vatten här.
		-- Sally Forth

%
Forskarna vet fortfarande mindre om vad som lockar män än de gör omvad som lockar myggor."Vad varje kvinna bör veta om Män"
		-- Dr. Joyce Brothers,

%
Hon har alltid trott på det gamla ordspråket - lämna dem när du ser bra ut.
		-- Anita Loos, "Gentlemen Prefer Blondes"

%
Hon varit gift så många gånger hon fick ris varumärken över hennes ansikte.
		-- Tom Waits

%
Hon härstammar från en lång rad som hennes mamma lyssnade på.
		-- Gypsy Rose Lee

%
Hon kom just in, kastade runt här med mig för ett par år, haftsjälv, gav det en slags vacker kvalitet och vänster. Upphetsad några mänsålänge.medverkan i "The Avengers".
		-- Patrick Macnee, reminiscing on Diana Rigg's

%
Hon tyckte om honom; Han var en man med många kvaliteter, även om de flesta av dem var dålig.
		-- Patrick Macnee, reminiscing on Diana Rigg's

%
Hon missade en ovärderlig möjlighet att ge honom en blick som du kanhar hälls på en våffla ...
		-- Patrick Macnee, reminiscing on Diana Rigg's

%
Hon har lärt sig att säga saker med ögonen som andra slösa tid att sättai ord.
		-- Patrick Macnee, reminiscing on Diana Rigg's

%
Hon är så tuff att hon inte kommer att ta "ja" för ett svar.
		-- Patrick Macnee, reminiscing on Diana Rigg's

%
Hon är den typ av tjej som klättrade på stegen av framgång fel genom fel.
		-- Mae West

%
Så många vackra kvinnor och så lite tid.
		-- John Barrymore

%
Så många män; så lite tid.
		-- John Barrymore

%
Så många kvinnor; så lite nerv.
		-- John Barrymore

%
Så många kvinnor; så lite tid!
		-- John Barrymore

%
"Så du inte behöver, Cindy, men jag undrar om du kanskevill gå till någonstans, du vet, med mig, någon gång. ""Ja, jag kan tänka mig en hel del värre saker, David.""Fredag, då?""Varför inte, David, det kan även vara kul."
		-- Dating in Minnesota

%
Vissa män är levande bevis på att en kvinna kan ta ett skämt.
		-- Dating in Minnesota

%
Vissa äktenskap made in heaven - men så är åska och blixtar.
		-- Dating in Minnesota

%
Vissa män är alla rätt i deras ställe - om de bara visste de rätta ställena!
		-- Mae West

%
Vissa män är så intresserade av deras fruar fortsatta lycka som dehyra detektiver att ta reda på orsaken till det.
		-- Mae West

%
Vissa män är så macho de ska få dig gravid bara för att döda en kanin.
		-- Maureen Murphy

%
En del män känner att det enda de är skyldiga den kvinna som gifter demär ett agg.
		-- Helen Rowland

%
Några av oss blir de män som vi ville gifta.
		-- Gloria Steinem

%
Ibland en cigarr bara en cigarr.
		-- Sigmund Freud

%
Ibland när jag tänker på vad den där tjejen betyder för mig, det är allt jag kan göraför att inte tala om för henne.
		-- Andy Capp

%
Stanford kvinnor är ansvariga för framgången för många Stanford män:de ger dem "bara ytterligare ett skäl" att bo i och studera varje natt.
		-- Andy Capp

%
Ta mitt ord för det, kan dummaste kvinnan hantera en smart man, men detbehöver en mycket smart kvinna för att hantera en dåre.
		-- Kipling

%
Tehee quod hon, och clapte den wyndow till.
		-- Geoffrey Chaucer

%
Den kvinnan talar åtta språk och kan inte säga "nej" i någon av dem.
		-- Dorothy Parker

%
Fördelen med att vara ogift är att när man ser en vacker flicka enbehöver inte sörja över att ha en ful ett hem.
		-- Paul Leautaud, "Propos d'un jour"

%
Vrede en kvinna är den största ondskan som du kan hota dinfiender.
		-- Bonnard

%
Den genomsnittliga flickan skulle hellre ha skönhet än hjärnor eftersom hon vetatt den genomsnittliga människan kan se mycket bättre än han kan tänka.
		-- Ladies' Home Journal

%
Den genomsnittliga kvinnan måste oundvikligen se hennes verkliga make med en vissförakt; han är allt annat än hennes ideal. Följaktligen kan hon inte hjälpakänslan av att hennes barn är grymt handikappad av det faktum att han ärderas far.
		-- H. L. Mencken

%
Den bästa mannen för jobbet är ofta en kvinna.
		-- H. L. Mencken

%
Det bästa med att vara skallig är, att när oväntade företaget anländer,Allt du behöver göra är att räta ut slips.
		-- H. L. Mencken

%
Den stora frågan är varför under evolutionen hanarna tillåtssig vara så helt skuggan av honorna. Varför de tolereradenna totala underkastelse, denna eländiga existens som utstötta som ärhungrig hela tiden?
		-- H. L. Mencken

%
Kedjorna äktenskap är så tung att det krävs två för att bära dem, ochibland tre.
		-- Alexandre Dumas

%
Dagarna strax före äktenskapet är som en kvick introduktion till entråkiga bok.
		-- Alexandre Dumas

%
Försvaret advokat hamrade bort på käranden:"Ni påstår," han hånade, "att min klient kom på dig med en trasig flaskai handen. Men är det inte sant, att du hade något i handen? ""Ja", mannen erkände, "sin fru. Mycket charmig, naturligtvis,men inte mycket bra i en kamp. "
		-- Alexandre Dumas

%
Skillnaden mellan laglig separation och skilsmässa är den juridiskaseparation ger man tid att gömma sina pengar.
		-- Alexandre Dumas

%
Varaktigheten av passion är proportionerlig med den ursprungliga motståndav kvinnan.
		-- Honor'e DeBalzac

%
Den eviga feminina drar oss uppåt.
		-- Goethe

%
Den första äktenskap är en triumf för fantasin över intelligens,och den andra är hoppets triumf över erfarenheten.
		-- Goethe

%
Herrarna såg varandra över med mikroskopisk slarv.
		-- Goethe

%
Flickan som minns sin första kyss nu har en dotter som inte ensminns sin första make.
		-- Goethe

%
Flickan som lutar sig att erövra vanligtvis bär en urringade klänning.
		-- Goethe

%
Flickan som svär ingen har någonsin älskat henne har en rätt att svära.
		-- Sophia Loren

%
Gudarna gav man eld och han uppfann brandbilar. De gav honomkärlek och han uppfann äktenskapet.
		-- Sophia Loren

%
Den lyckligaste tiden av en människas liv är efter hans första skilsmässa.
		-- J. K. Galbraith

%
Den tyngsta objekt i världen är kroppen av kvinnan du har upphörtatt älska.
		-- Marquis de Lac de Clapiers Vauvenargues

%
Smekmånaden är faktiskt inte över förrän vi upphör att kväva våra suckaroch börja att kväva våra gäspningar.
		-- Helen Rowland

%
Smekmånaden är över när han telefoner för att säga att han kommer för sent till kvällsmat ochHon har redan lämnat en anteckning om att det är i kylskåpet.
		-- Bill Lawrence

%
Mannen som inte berätta för sin fru allt förmodligen skäl somVad hon inte vet kommer inte att skada honom.
		-- Leo J. Burke

%
Den lilla flickan förväntar sig ingen försäkran om ömhet från sin docka.Hon älskar det - och det är allt. Det är därför som vi skulle älska.
		-- DeGourmont

%
Majoriteten av män påminner mig om en orangutang försöker spela fiol.
		-- Honor'e DeBalzac

%
Mannen som förstår en kvinna är kvalificerad att förstå ganska braallt.
		-- Yeats

%
Den mogna bohemiska är ett vars kvinna arbetar heltid.
		-- Yeats

%
Den vanligaste formen av frieri: "DU VAD !?"
		-- Yeats

%
Den mest farliga livsmedel är bröllopstårta.
		-- American proverb

%
De svåraste åren av äktenskap är de efter bröllopet.
		-- American proverb

%
Den mest lyckligt äktenskap jag kan tänka mig att själv skulle vara förbundetav en döv man till en blind kvinna.
		-- Samuel Taylor Coleridge

%
Det viktigaste i en relation mellan en man och en kvinnaär att en av dem vara bra på att ta order.
		-- Linda Festa

%
De mest populära arbetsbesparande enhet idag är fortfarande en man med pengar.
		-- Joey Adams, "Cindy and I"

%
Modern av året bör vara en steriliserad kvinna med två adopterade barn.
		-- Paul Ehrlich

%
Den charm äktenskapet är att det gör ett liv av bedrägeri en nödvändighet.
		-- Oscar Wilde

%
Den enda verkliga argument för äktenskapet är att det fortfarande den bästa metodenför att bekanta.
		-- Heywood Broun

%
Den enda riktigt mäster buller en man gör i ett hus är bullretav sin nyckel, när han är fortfarande på landning, trevande för låset.
		-- Colette

%
Den perfekta människan är den sanna partnern. Inte en säng partner eller en rolig partner,men en man som kommer att axla bördan lika med [du] och har somkvalitet av glädje.
		-- Erica Jong

%
Den person som gifter sig för pengar tjänar vanligtvis vartenda öre av det.
		-- Erica Jong

%
De vackraste kvinnor är nästan alltid det tråkigaste, och det är därförvissa människor känner att det finns ingen Gud.
		-- Woody Allen, "Without Feathers"

%
Den Ruffed Pandanga av Borneo och Rotherham breder ut sina fjädrar ihans uppvaktning dans och imiterar Winston Churchill och Tommy Cooperena benet. Den padanga dör ut eftersom den kvinnliga padanga inteta det för allvarligt.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
De sex stora gåvor en irländsk flicka är skönhet, mjuk röst, söt tal,visdom, handarbete, och kyskhet.
		-- Theodore Roosevelt, 1907

%
Det säkraste tecknet på att en man är kär är när han skiljer sig från sin fru.
		-- Theodore Roosevelt, 1907

%
Problemet med vissa kvinnor är att de får alla glada om ingenting- Och sedan gifta sig med honom.
		-- Cher

%
Sanningen om en kvinna varar ofta längre än kvinnan är sant.
		-- Cher

%
De två saker som kan få dig i trubbel snabbare än något annatär snabba kvinnor och långsamma hästar.
		-- Cher

%
Sättet att bekämpa en kvinna är med din hatt. Ta det och köra.
		-- Cher

%
Kvinnan du köper - och hon är den billigaste - tar en stordel pengar. Kvinnan som ger sig tar all din tid.
		-- Balzac

%
Det finns några saker som aldrig går ur stil, och en kvinnlig kvinnaär en av dem.
		-- Ralston

%
Det finns fyra steg till ett äktenskap. Först finns det affären, så finns detäktenskapet, då barn och slutligen den fjärde etappen, utan som dukan inte känna en kvinna, skilsmässa.
		-- Norman Mailer

%
Det finns tre saker som jag har alltid älskat och aldrig förstått -konst, musik och kvinnor.
		-- Norman Mailer

%
Det finns tre saker män kan göra med kvinnor: älska dem, lida för dem,eller förvandla dem till litteratur.
		-- Stephen Stills

%
Det finns två tillfällen då man inte förstår en kvinna - innanäktenskap och efter äktenskapet.
		-- Stephen Stills

%
Det går bra tid som var hade alla.
		-- Bette Davis, remarking on a passing starlet

%
Det finns en stor skillnad mellan den vilda och civiliserade människan, men detär aldrig klart för sina fruar förrän efter frukost.
		-- Helen Rowland

%
Det finns ingen realiserbara kraft som människan kan inte, i tid, mode verktygenatt uppnå, eller någon makt så säkra att blotta apan inte kommer att missbruka det.Så det står skrivet i de genetiska kort - bara fysik och krig hålla honom ikolla upp. Och även fru som vill ha honom hem med fem, naturligtvis.
		-- Encyclopadia Apocryphia, 1990 ed.

%
Det finns inget sådant som en ful kvinna - det finns bara de som görinte vet hur man gör sig attraktiv.
		-- Christian Dior

%
Det finns inte mycket att välja mellan en kvinna som lurar oss för en annan,och en kvinna som lurar en annan för oss själva.
		-- Augier

%
Det finns bara ett sätt att trösta en änka. Men kom ihåg risken.
		-- Robert Heinlein

%
Det finns inget som en flicka med en djup urringning att hålla en man på tårna.
		-- Robert Heinlein

%
Det finns inget som en god dos av en annan kvinna att göra en människa att uppskattahans fru.
		-- Clare Booth Luce

%
Det finns inget som god mat, gott vin och en dålig flicka.
		-- Clare Booth Luce

%
Det finns en tröst om äktenskap. När du tittar runt du kanalltid se någon som gjorde värre.
		-- Warren H. Goldsmith

%
Det finns en dåre åtminstone i varje gift par.
		-- Warren H. Goldsmith

%
Det finns bara ett sätt att få ett lyckligt äktenskap och så fort jag läravad det är jag ska gifta igen.
		-- Clint Eastwood

%
Det finns för mycket skönhet på denna jord för ensamma män att bära.
		-- Richard Le Gallienne

%
Den här killen går in i hans hus och skriker till sin fru, "Kathy, packa upp dinväskor! Jag vann bara Kalifornien lotteri! ""Älskling!", Kathy utropar, "Ska jag packa för varmt väder eller kallt?""Jag bryr mig inte", svarar mannen. "Bara så länge som du är uteav huset med middag! "
		-- Richard Le Gallienne

%
'Tis saligare att ge än få, till exempel, presenterar bröllop.
		-- H. L. Mencken

%
Att vara vacker är nog! om en kvinna kan göra det bra som borde krävamer från henne? Du vill inte en ros att sjunga.
		-- Thackeray

%
För att betraktas som framgångsrik, måste en kvinna vara mycket bättre på sitt jobbän en man skulle behöva vara. Lyckligtvis är detta inte svårt.
		-- Thackeray

%
För att bli framgångsrik, har en kvinna att vara mycket bättre på sitt jobb än en människa.
		-- Golda Meir

%
Att fela är mänskligt - men det känns gudomligt.
		-- Mae West

%
Att ta reda på en flicka fel, beröm henne till hennes väninnor.
		-- Benjamin Franklin

%
För många är total avhållsamhet lättare än perfekt måtta.
		-- St. Augustine

%
Till våra älsklingar och hustrur. Kan de träffas aldrig.
		-- 19th century toast

%
Idag när en man gifter sig får han ett hem, en hushållerska, en kock, en jublandetrupp och en annan lönecheck. När en kvinna gifter sig, får hon en boarder.
		-- 19th century toast

%
För mycket av det goda är underbart.
		-- Mae West

%
Lita på din make, älska din man, och få så mycket som möjligt ieget namn.
		-- Joan Rivers

%
Tjugo år av romantik göra en kvinna ser ut som en ruin; men tjugo år aväktenskap göra henne något som en offentlig byggnad.
		-- Oscar Wilde

%
Två säker sätt att berätta en riktigt sexig man; det första är, han har ett dåligt minne.Jag glömmer den andra.
		-- Oscar Wilde

%
Fram till Eva kom, var detta en mans värld.
		-- Richard Armour

%
Valerie: AWW, Tom, du kommer maudlin på mig ...Tom: Jag förbehåller oss rätten att vaxa maudlin som jag avta vältalig ...
		-- Tom Chapin

%
Mycket få moderna kvinnor antingen gillar eller önskan äktenskap, särskilt efterceremoni har utförts. Främst kvinnor önskar uppmärksamhet och tillgivenhet.Äktenskapet är något de accepterar när det inte finns något alternativ. Verkligen,det är ett slöseri med tid, och farligt, att gifta dem. Det lämnar en öppentill en rival. Män, bra eller dåliga, alltid har rivaler. Älskare, aldrig.
		-- Helen Lawrenson, "Esquire"

%
Vi var lyckligt gifta i åtta månader. Tyvärr var vi giftaför fyra och ett halvt år.
		-- Nick Faldo

%
Vi är alla söker en kvinna som kan sitta i en minikjol och pratafilosofi, verkställande både med tillförsikt och stil.
		-- Nick Faldo

%
Bröllop är öde, och hänger på samma sätt.
		-- John Heywood

%
Vigselringar är världens minsta handbojor.
		-- John Heywood

%
Tja, det är svårt för en vanlig människa att tro att kvinnan inte har lika rättigheter.
		-- Dwight D. Eisenhower

%
Vad en olycka att vara en kvinna! Och ändå är det värsta olycka inteförstå vad en olycka det är.
		-- Kierkegaard, 1813-1855.

%
Vad ger du en man som har allt? Penicillin.
		-- Jerry Lester

%
"Vad ger du en man som har allt?" den vackra tonåringfrågade sin mamma."Uppmuntran, kära", svarade hon.
		-- Jerry Lester

%
Vilka dumheter människor talar om lyckliga äktenskap! En man kan vara nöjd meden kvinna så länge han inte älskar henne.
		-- Oscar Wilde

%
Vad passerar för kvinna intuition är ofta ingenting mer än människansgenomskinlighet.
		-- George Nathan

%
Vad förlag letar efter dessa dagar är inte radikal feminism. Desscorporate feminism - ett varumärke av feminismen som syftar till att sälja böcker ochtidskrifter, tredelade kostymer, flygbiljetter, Scotch, cigaretter och,viktigast, corporate America budskap, som lyder: Ja, kvinnordiskrimineras i det förflutna, men det olyckligt misstag har varitåtgärdas; nu varje kvinna kan uppnå rikedom, prestige och makt genom dintindividuell snarare än kollektiv insats.
		-- Susan Gordon

%
Oavsett kvinnor gör de måste göra dubbelt så bra som män att ses halvlika bra. Lyckligtvis är detta inte svårt.
		-- Charlotte Whitton

%
När en flicka kan läsa handstil på väggen, kan hon vara i felvilorum.
		-- Charlotte Whitton

%
När en flicka gifter hon byter uppmärksamhet av många män förinattentions av en.
		-- Helen Rowland

%
När en man stjäl din fru, det finns inget bättre hämnd än att låta honomhålla henne.
		-- Sacha Guitry

%
När en kvinna ger mig en present jag har alltid två överraskningar:första är närvarande, och efteråt, att behöva betala för det.
		-- Donnay

%
När en kvinna gifter sig igen beror det på att hon avskydde sin första make.När en man gifter sig igen, är det för att han älskade sin första hustru.
		-- Oscar Wilde

%
När du väljer mellan två onda ting, jag gillar alltid att ta en jag har aldrigförsökt innan.
		-- Mae West, "Klondike Annie"

%
När Gud skapade två könen, kan han ha varit överdriven det.
		-- Charles Merrill Smith

%
När Gud såg hur felaktig var man Han försökte igen och gjorde kvinnan. attvarför han då slutade det finns två åsikter. En av dem är kvinnans.
		-- DeGourmont

%
När jag var en ung man, lovade jag att aldrig gifta tills jag hittade den perfektakvinna. Tja, jag hittade henne - men tyvärr, hon väntade på den perfekta mannen.
		-- Robert Schuman

%
När jag är bra, jag är bra; men när jag är dålig, jag är bättre.
		-- Mae West

%
När det gäller trasiga äktenskap flesta män kommer att dela skulden -halv hans fru fel, och halv hennes mors.
		-- Mae West

%
När Äktenskapet kriminaliseras, kommer bara Outlaws har inlaws.
		-- Mae West

%
När mitt första rumskamrat vid Cornell fick veta att jag var jude, var hon påhennes begäran, flyttade till ett annat rum. Hon berättade att hon trodde inte att honhade någonsin sett en Judisk innan. Min enda svar var att börja bära enliten davidsstjärna på en kedja runt halsen. Jag hade inte blivit en merobservera Judisk; snarare, upptäcker att märkningen av Judisk var kränkande förandra fick mig att vilja låta folk veta vem jag var och vad jag trodde på.På samma sätt, efter att ha talat med dessa unga kvinnor - varav berättade attHon trodde inte att hon någonsin hade träffat en feminist - jag har tagit till att identifierasjälv som feminist i de mest osannolika situationer.
		-- Susan Bolotin, "Voices From the Post-Feminist Generation"

%
När man vet kvinnor en ömhet män, men när man studerar män,en ursäkter kvinnor.
		-- Horne Tooke

%
När ljusen är ute alla kvinnor är rättvist.
		-- Plutarch

%
När saleman bil sönder, gick han till närmaste hus för att frågaom han kunde stanna natten. Bonden kom överens om att sätta upp honom. "Jag bor ensam,"fortsatte han, "du kan ha sovrum på toppen av trappan, tillhöger.""Åh, strunt", den besviken försäljaren sa. "Jag tror jag ärfel skämt. "
		-- Plutarch

%
När det finns en gammal fröken i huset, är en vakthund onödig.
		-- Balzac

%
När två personer är under inflytande av de mest våldsamma, mest galen,mest bedrägliga, och mest övergående av passioner, är de skyldiga att sväraatt de kommer att förbli i det glada, onormal, och ansträngande tillståndkontinuerligt tills döden skiljer dem del.
		-- George Bernard Shaw

%
När kvinnor kysser det alltid påminner en av pris kämpar skakar hand.
		-- H. L. Mencken, "Sententiae"

%
När kvinnor älskar oss, de förlåter oss allt, även våra brott; när de görinte älska oss, de ger oss kredit för ingenting, inte ens våra dygder.
		-- Honor'e de Balzac

%
När du är uttråkad med dig själv, att gifta sig, och bli uttråkad med någon annan.
		-- David Pryce-Jones

%
När du är gift med någon, de tar dig för givet ... närdu lever med någon det är fantastiskt ... de är så räddaatt förlora dig de har att hålla dig nöjd hela tiden.
		-- Nell Dunn, "Poor Cow"

%
När jag går en kille, tror jag, är detta den man jag vill att mina barnatt tillbringa sina helger med?
		-- Rita Rudner

%
Var är mannen kan underlätta ett hjärta som en satängkappa?
		-- Dorothy Parker, "The Satin Dress"

%
Varför man vill ha en fru är ett stort mysterium för vissa människor. Varför en manvill * ___ två * fruar är en bigamystery.
		-- Dorothy Parker, "The Satin Dress"

%
Varför finns det inte några billiga och enkelt sätt att bevisa hur mycket hon betyder för mig?
		-- Dorothy Parker, "The Satin Dress"

%
Varför vill du inte låta mig kyssa dig godnatt? Är det något som jag sade?
		-- Tom Ryan

%
Med slutet av fotbollssäsongen, en stjärnspelare för college lagetfirade uppmjukning av laget utegångsförbud genom att delta i en sena campuspart. Strax efter ankomsten, blev han fångade av en vacker coed ochlättade i en konversation med henne genom att fråga om hon träffade många datum påparter."Åh, jag har en tre punkt åtta, så jag är mycket mer lockas tillstarka akademiska typer än de dumma parti djur ", sade hon." Vad ärdin G.P.A.? "Grina öra till öra, skröt Jock, "Jag får ungefär tjugofem istaden och fyrtio på motorvägen. "
		-- Tom Ryan

%
Kvinna inspirerar oss till stora saker, och hindrar oss från att nå dem.
		-- Dumas

%
Kvinnan var Guds andra misstag.
		-- Nietzsche

%
Kvinnan togs ut av människan - inte ut ur hans huvud, att härska över honom; inte hellerav hans fötter, att trampas under av honom; men ur hans sida, att varalika med honom - under armen, att han skulle skydda henne, och nära hans hjärtaatt han skulle älska henne.
		-- Henry

%
Kvinnans råd har ringa värde, men den som inte tar det är en dåre.
		-- Cervantes

%
Kvinnor är alla lika. När de är pigor de är mild som mjölk: en gång göra demfruar, och de lutar ryggen mot sina äktenskapscertifikat, ochtrotsa dig.
		-- Jerrold

%
Kvinnor är alltid angelägna om att uppmana ungkarlar till äktenskap; är det från välgörenhet,eller hämnd?
		-- Gustave Vapereau

%
Kvinnor är precis som män, endast annorlunda.
		-- Gustave Vapereau

%
Kvinnor är som elefanter till mig: Jag gillar att titta på dem, men jag skulle intevill äga en.
		-- W. C. Fields

%
Kvinnor är inte mycket, men de är de bästa motsatta könet vi har.
		-- Herold

%
Kvinnor är klokare än män eftersom de vet mindre och förstå mer.
		-- Stephens

%
Kvinnor är inte så ren som de brukade vara.
		-- Pogo

%
Kvinnor kan hålla en hemlighet lika bra som män, men det krävs mer av dematt göra det.
		-- Pogo

%
Kvinnor klagar sex mer än män. Deras gnäller falla i tvåkategorier: (1) Inte tillräckligt och (2) För mycket.
		-- Ann Landers

%
Kvinnor ger sig till Gud när Djävulen vill inget mer att göra med dem.
		-- Arnould

%
Kvinnor ge män själva guldet av deras liv. Eventuellt; men dealltid vill ha tillbaka så mycket liten förändring.
		-- Oscar Wilde

%
Kvinnor i kärlek består av en liten suckande, lite gråt, lite döende- Och en hel del att ligga.
		-- Ansey

%
Kvinnor resonera med hjärtat och är mycket mindre ofta fel än män somresonera med huvudet.
		-- DeLescure

%
Kvinnor förlåta ibland en man som tvingar möjlighet, men aldrig en människasom missar ett.
		-- Charles De Talleyrand-Perigord

%
Kvinnor behandla oss lika mänskligheten behandlar sina gudar. De dyrkar oss och äralltid stör oss att göra något för dem.
		-- Oscar Wilde

%
Kvinnor vill att deras män att vara poliser. De vill att du ska straffa dem och berättadem vad gränserna går. Det enda som kvinnor hatar värre från en människaän bli slagen är när du får på knä och säga att du är ledsen.
		-- Mort Sahl

%
Kvinnor avfall mäns liv och tror att de har ersätts dem med ett fåtalnådens ord.
		-- Honor'e de Balzac

%
Kvinnor som vill vara lika med män saknar fantasi.
		-- Honor'e de Balzac

%
Kvinnor vill bli älskad utan varför eller varför; inte för att de ärsöt, eller bra, eller belevad, eller graciös, eller intelligent, men eftersomde själva.
		-- Amiel

%
Kvinnors dygd är människans största uppfinning.
		-- Cornelia Otis Skinner

%
Kvinnor, lurade av män, vill gifta sig med dem; det är ett slags hämndså gott som alla andra.
		-- Philippe De Remi

%
Kvinnor, när de inte är kär, har alla kallblodigt av en erfarenadvokat.
		-- Honor'e de Balzac

%
Kvinnor, när de har gjort ett får av en man, alltid tala om för honom att han är enlejon med en vilja av järn.
		-- Honor'e de Balzac

%
	"Du är så underbar.""Ja.""Ja! Och du tar en komplimang, alltför! Jag gillar det i en gudinna."
		-- Honor'e de Balzac

%
Det är inte tillåtet att döda en kvinna som har kränkt dig, men ingentingförbjuder dig att reflektera att hon växer äldre varje minut. Du ärhämnd fjorton hundra fyrtio gånger om dagen.
		-- Ambrose Bierce

%
Du frågar vad en trevlig tjej kommer att göra? Hon kommer inte att ge en tum, men hon kommer intesäger nej.
		-- Marcus Valerius Martialis

%
Du kan ha en hund som en vän. Du kan ha whisky som en vän. MenOm du har en kvinna som en vän, du kommer att hamna berusad och kyssasdin hund.
		-- foolin' around

%
Du kan aldrig lita på en kvinna; hon kan vara sant för dig.
		-- foolin' around

%
Du kan inte kyssa en flicka oväntat - endast tidigare än hon trodde att du skulle.
		-- foolin' around

%
Du behöver bara mumla några ord i kyrkan för att gifta och några ordi sömnen för att få frånskild.
		-- foolin' around

%
Du vet precis när en relation är på väg att ta slut. Min flickvän ringde migpå jobbet och frågade mig hur man byta en glödlampa i badrummet. "Det är väldigtenkel, "sa jag." Du börjar med att fylla upp badkaret med vatten ... "
		-- foolin' around

%
Du vet vad vi kan vara som: Se en kille och tycker att han är söt en minut,nästa minut våra hjärnor har vi gift med barn, följande minuten vi serhan har ett utomäktenskapligt förhållande. Genom säger gång någon "Jag skulle vilja att niMöt Cecil, "vi ropa:" Du är sen igen med barnet stöd! "
		-- Cynthia Heimel, "A Girl's Guide to Chaos"

%
Du vet att du får gammal när du är pappa, och du mäter din dotterför läger kläder, och det finns vissa mätningar bara hennes mor är tillåtetatt ta.
		-- Cynthia Heimel, "A Girl's Guide to Chaos"

%
Du vet, naturligtvis, att Tasmanians, som aldrig begått äktenskapsbrott,är nu utdöda.
		-- M. Somerset Maugham

%
Du bodde med en man som bar vitbälten? Laura, jag är besviken på dig.
		-- Remington Steele

%
Du tror Oidipus hade ett problem - Adam var Evas mamma.
		-- Remington Steele

%
"Du är just den typ av person som jag föreställt gifta, när jag var liten ...utom, du vet, inte grönt ... och utan alla fläckar av svamp. "
		-- Swamp Thing

%
Unga män och unga kvinnor kan arbeta systematiskt sex dagar ivecka och stiga färskt på morgonen, men låt dem delta moderna danser förbara några timmar varje kväll och se vad som händer. Vals, polka,Galopp och andra danser av samma slag kommer att bli katastrofala i deras effektertill båda könen. Hälsa och vigör kommer att försvinna som dagg innan solen.Det är inte ovanligt övning som skadar dansaren, mensnarare kommer i nära kontakt med det motsatta könet. Det ärraseri lust sugen oavbrutet för mer glädje som undergräversjäl, kropp, senor och nerver. Erfarenhet och statistik visarbortom allt tvivel att passionerade alltför dansande flickor knappast kan nåtjugofem år och män trettio-en. Även om de kom attålder kommer de i de flesta fall brytas hälsa fysiskt och moraliskt.Detta är påståendet framstående läkare i detta land.
		-- Quote from a 1910 periodical

%
Unga män vill vara trogna och är inte; gamla män vill vara trolös ochkan inte.
		-- Oscar Wilde

%
Ungdom hade varit en vana av hennes så länge att hon kunde inte del med det.
		-- Oscar Wilde

%
