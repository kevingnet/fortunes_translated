En bank är en kollega som lånar du hans paraply när solen skineroch vill ha tillbaka den minut det börjar regna.
		-- Mark Twain

%
En klassiker är något som alla vill ha lästoch ingen vill läsa.
		-- Mark Twain, "The Disappearance of Literature"

%
En häst! En häst! Mitt kungarike för en häst!
		-- Wm. Shakespeare, "Richard III"

%
Hundra år från nu är det mycket troligt att [av Twain verk] "TheJumping Frog "enbart kommer att bli ihågkommen.
		-- Harry Thurston Peck (Editor of "The Bookman"), January 1901.

%
A är för Apple.
		-- Hester Pryne

%
Ett slags Batman samtida bokstäver.
		-- Philip Larkin on Anthony Burgess

%
En lätt hustru bliver en tung make.
		-- Wm. Shakespeare, "The Merchant of Venice"

%
En man läste The Canterbury Tales en lördag morgon, när hansfru frågade "Vad har du där?" Svarade han, "Just my cup och Chaucer."
		-- Wm. Shakespeare, "The Merchant of Venice"

%
... En högtidlig, unsmiling, skenheliga gamla isberg som såg ut som om hanväntade på en ledig plats i treenigheten.
		-- Mark Twain

%
Två städer LITE (tm)- Vid Charles DickensEn advokat som ser ut som en fransk adelsman utförs i hans ställe.Förvandlingen LITE (tm)- Av Franz KafkaEn man förvandlas till en bugg och hans familj blir irriterad.Sagan om Ringen LITE (tm)- Av J. R. R. TolkienVissa killar ta en lång semester för att kasta en ring i en vulkan.Hamlet LITE (tm)- Av Wm. ShakespeareEn högskolestudent på semester med familjeproblem, en screwyflickvän och en mor som inte kommer att agera hennes ålder.
		-- Mark Twain

%
Två städer LITE (tm)- Vid Charles DickensEn man kär i en tjej som älskar en annan man som ser ut precissom han har huvudet avhuggna i Frankrike på grund av en genomsnittligdam som stickar.Brott och straff LITE (tm)- Vid Fyodor DostoevskiEn man skickar en otäck brev till en pantbank, men senarekänns skyldig och ber om ursäkt.Odyssey LITE (tm)- Av HomerEfter att ha arbetat sent, blir en tapper krigare förlorade på väg hem.
		-- Mark Twain

%
När allt kommer omkring, allt han gjorde var sträng tillsammans en hel del gamla, välkända citat.
		-- H. L. Mencken, on Shakespeare

%
Ack, hur kärleken kan leka med sig själv!
		-- William Shakespeare, "The Two Gentlemen of Verona"

%
Alla generaliseringar är falska, inklusive denna.
		-- Mark Twain

%
Allt jag vet är vad orden vet, och döda ting, och attgör en vacker liten summa, med en början och ett mellersta ochett slut, som i den välbyggda fras och lång sonaten av de döda.
		-- Samuel Beckett

%
Alla säger, "Hur svårt det är att vi måste dö" - en konstig klagomål komma frånmunnen från personer som har varit tvungna att leva.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
"... Alla moderna olägenheter ..."
		-- Mark Twain

%
Allt som är med mer ande jagade än haft.
		-- Shakespeare, "Merchant of Venice"

%
gör alltid rätt. Detta kommer att tillfredsställa vissa människor och förvåna resten.
		-- Mark Twain

%
Alltid slöhet av dåren är brynet av förstånd.
		-- William Shakespeare, "As You Like It"

%
"... En erfaren, flitig, ambitiös, och ofta ganska oftapittoreska lögnare. "
		-- Mark Twain

%
En ärlig berättelse hastigheter bäst att tydligt höra.
		-- William Shakespeare, "Henry VI"

%
Och tror ni (FOP som jag) att jag kunde vara Scarlet pumpernickel?
		-- William Shakespeare, "Henry VI"

%
Alla som har haft en tjur i svansen vet fem eller sex fler sakerän någon som inte har.
		-- Mark Twain

%
april 1Detta är den dag då vi påminns om vad vi är på de andra trehundra och sextiofyra.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Som flyger till hänsynslösa pojkar är vi till gudarna; de dödar oss för sin sport.
		-- Shakespeare, "King Lear"

%
När det gäller Adjektiv: när du är osäker, slå ut.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
På en gång slog det mig vilken kvalitet gick att bilda en man av prestation,särskilt i litteraturen, och som Shakespeare hade så enormt- Jag menar negativ kapacitet, det vill säga när en man är i stånd atti osäkerhet, mysterier, tvivel, utan någon irriterad nårefter fakta och förnuft.
		-- John Keats

%
VAKEN! RÄDSLA! BRAND! Fiender! VAKEN!FEAR! BRAND! Fiender!VAKNA! VAKEN!
		-- J. R. R. Tolkien

%
Awash med ofokuserad önskan, Everett vred loben av hans enda kvarvarandeörat och kände närvaron av någon annan bakom honom, vilket orsakade skräckatt driva igenom sitt nervsystem som en störtflod dånande nermid-gaffel av Feather River innan slutförandet av Oroville Dam1959.dålig fiction tävling.
		-- Grand Panjandrum's Special Award, 1984 Bulwer-Lytton

%
Var försiktig med att läsa hälsa böcker, kan du dö av ett tryckfel.
		-- Mark Twain

%
Se, dåren säger, "Sätt inte alla dina ägg i en korg" - som ärmen ett sätt att säga, "Scatter dina pengar och din uppmärksamhet;" men den viseman säger, "lägga alla ägg i en korg och - titta på det BASKET."
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Stor bok, stora hål.
		-- Callimachus

%
Men för min egen del, var det grekiska för mig.
		-- William Shakespeare, "Julius Caesar"

%
Genom att försöka kan vi enkelt lära sig att uthärda motgångar. En annan mans, menar jag.
		-- Mark Twain

%
Civilisation är den obegränsade multiplikation onödiga nödvändigheter.
		-- Mark Twain

%
Kläderna gör mannen. Nakna människor har liten eller ingen inverkan på samhället.
		-- Mark Twain

%
Kondensera soppa, inte böcker!
		-- Mark Twain

%
Samvetet bliver fegisar av oss alla.
		-- Shakespeare

%
Överväga väl proportionerna av saker. Det är bättre att vara en ung juni-bugän en gammal fågel av paradiset.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Mod är motstånd att frukta, behärskningen av rädsla - inte avsaknaden av rädsla. utom envarelse vara del feg det är inte en komplimang att säga att det är modig; det är endasten lös missbruk av ordet. Tänk på lopp - ojämförligtmodigaste av alla varelser av Gud, om okunnighet om rädsla var mod.Oavsett om du sover eller vaken han kommer att attackera dig, att bry sig ingenting för det faktumatt i bulk och styrka du är till honom som är hopade arméer på jordentill en sugande barn; han bor både dag och natt och alla dagar och nätter imycket varvet av fara och den omedelbara närvaron av döden, och ändå är inte merrädd än vad man som vandrar på gatorna i en stad som hotas aven jordbävning tio århundraden före. När vi talar om Clive, Nelson, och Putnamsom män som "inte vet vad rädsla var," vi borde alltid att lägga loppan - ochsatte honom i spetsen för processionen.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Fördröjning inte, Caesar. Läs den direkt.Här är ett brev, läsa den på din fritid.[Citerat i "VMS interna och datastrukturer", V4.4, närmed hänvisning till I / O-systemtjänster.]
		-- Shakespeare, "Merchant of Venice" 5,1

%
Delores seglade längs ytan av sitt liv som en flat sten för evigthoppa längs slät vatten, porlande verkligheten sporadiskt men omedvetnadet konsekvent, tills hon slutligen förlorade fart, sjönk, och på grund av enöverdos av flouride som barn som fick henne att lida av kroniskapati, dömd sig ligga alltid på golvet i hennes liv som värdelössom en bilaga och som ensam som en femhundra pund skivstång i ensteroid-gratis gym.
		-- Winning sentence, 1990 Bulwer-Lytton bad fiction contest.

%
Inte gå omkring och säga att världen är skyldig dig en levande. Världen är skyldig digingenting. Det var här först.
		-- Mark Twain

%
"Älvor och drakar!" Jag säger till honom. "Kål och potatis är bättreför dig och mig. "
		-- J. R. R. Tolkien

%
Engelsk litteratur är att utföra loppa.
		-- Sean O'Casey on P. G. Wodehouse

%
Även det tydligaste och mest perfekta indicier är sannolikt att vara påfel, trots allt, och därför borde tas emot med stor försiktighet. TaVid varje penna, slipas av någon kvinna; om du har vittnen, kommer duhitta hon gjorde det med en kniv, men om du tar helt enkelt den del av pennan,ni kommer att säga att hon gjorde det med tänderna.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Varje moln alstrar inte en storm.
		-- William Shakespeare, "Henry VI"

%
Varje varför har en varför.
		-- William Shakespeare, "A Comedy of Errors"

%
Extrem rädsla kan varken slåss eller fly.
		-- William Shakespeare, "The Rape of Lucrece"

%
F.S. Fitzgerald till Hemingway:"Ernest, de rika skiljer sig från oss."Hemingway:"Ja. De har mer pengar."
		-- William Shakespeare, "The Rape of Lucrece"

%
Fame är en ånga; popularitet en olycka; det enda jordiska säkerhet ärglömska.
		-- Mark Twain

%
Förtrogenhet föder förakt - och barn.
		-- Mark Twain

%
Få saker är svårare att stå ut med än irritation av ett bra exempel.
		-- "Mark Twain, Pudd'nhead Wilson's Calendar"

%
För en lätt hjärta lever länge.
		-- Shakespeare, "Love's Labour's Lost"

%
För mod mounteth med tillfälle.
		-- William Shakespeare, "King John"

%
För mode Minas Tirith var sådan att det byggdes på sju nivåer,varje grävde i en kulle, och om varje sattes en vägg, och i varje väggvar en grind.[Citerat i "VMS interna och datastrukturer", V4.4, närmed hänvisning till systemöversikt.]
		-- J.R.R. Tolkien, "The Return of the King"

%
För det finns stunder då man kan varken tänka eller känna. Och om man kanvarken tänka eller känna, hon tänkte, där är en?[Citerat i "VMS interna och datastrukturer", V4.4, närhänvisning till kraftfel återhämtning.]
		-- Virginia Woolf, "To the Lighthouse"

%
För år en hemlig skam förstörde min peace--Jag skulle inte läsa Eliot, Auden eller MacNiece.Men nu tror jag en tanke som ger mig hopp:Inte heller hade Chaucer, Shakespeare, Milton, Pope.
		-- Justin Richardson.

%
Gå inte till älvorna för råd, för de kommer att säga både ja och nej.
		-- J.R.R. Tolkien

%
Borta med vinden LITE (tm)- Av Margaret MitchellEn kvinna gillar bara män hon kan inte ha och södra blir skrotade.Gåva av Magi LITE (tm)- O. HenryEn man och hustru glömt att registrera sina gåva preferenser.Den gamle och havet LITE (tm)- Ernest HemingwayEn gammal man går fiske, men har inte mycket tur.
		-- J.R.R. Tolkien

%
Tacksamhet och förräderi är bara de två ändarna av samma processionen.Ni har sett allt det som är värt att stanna när bandet och pråligatjänstemän har gått.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Sorg kan ta hand om sig själv; men för att få det fulla värdet av en glädje som du måstehar någon att dela den med.
		-- Mark Twain

%
Vana är vana, och inte kastas ut genom fönstret av någon människa, men lirkadened-trappor ett steg i taget.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar

%
Hain't vi fick alla dårar i stan på vår sida? Och hain't att en stortillräckligt majoritet i någon stad?
		-- Mark Twain, "Huckleberry Finn"

%
Harpa inte på den strängen.
		-- William Shakespeare, "Henry VI"

%
Har en plats för allt och hålla sak någon annanstans; det här är interåd, är det bara sed.
		-- Mark Twain

%
Har ingenting, ingenting kan han förlora.
		-- William Shakespeare, "Henry VI"

%
Han drager ut tråden av hans informationsnivån finare än stapelvara i sinargument.
		-- William Shakespeare, "Love's Labour's Lost"

%
Han har ätit mig ut ur hus och hem.
		-- William Shakespeare, "Henry IV"

%
Han är nu stiger från rikedom till fattigdom.
		-- Mark Twain

%
Han skämt på ärr som aldrig kände ett sår.
		-- Shakespeare, "Romeo and Juliet, II. 2"

%
Han som bryter en sak att ta reda på vad det är har lämnat väg visdom.
		-- J.R.R. Tolkien

%
Han som är svindlande tror världen vänder.
		-- William Shakespeare, "The Taming of the Shrew"

%
Han var en del av min dröm, naturligtvis - men då var jag en del av hans dröm också.
		-- Lewis Carroll

%
Helvetet är tom och alla djävlar är här.
		-- Wm. Shakespeare, "The Tempest"

%
Hans anhängare kallade honom Mahasamatman och sa att han var en gud. han föredrogatt släppa Maha- och -atman dock och kallade sig Sam. han aldrigpåstod sig vara en gud. Men sedan, hävdade han aldrig inte vara en gud. omständig-ämnen var som den var, kunde ingen antagning vara till någon nytta.Tystnad, men kunde. Det var i dagarna av regn som sina bönergick upp, inte från finger av knotiga bön sladdar eller spinning avbön hjul, men från den stora be-maskin i klostret Ratri,gudinna av natten. högfrekventa böner de riktades uppåt genomatmosfären och bortom den, passerar in i den gyllene moln kallasBridge of the Gods, som cirklar hela världen, ses som en bronsregnbåge på natten och är den plats där den röda solen blir apelsin vid middagstid.Några av munkarna tvivlade ortodoxi denna bön teknik ...
		-- Roger Zelazny, "Lord of Light"

%
Hur apt de fattiga är att vara stolt.
		-- William Shakespeare, "Twelfth-Night"

%
Jag önskar att vi kan vara bättre främlingar.
		-- William Shakespeare, "As You Like It"

%
Jag vet inte hälften av er hälften så bra som jag skulle vilja; och jag gillar mindreän hälften av er hälften så bra som du förtjänar.
		-- J. R. R. Tolkien

%
Jag dote på hans mycket frånvaro.
		-- William Shakespeare, "The Merchant of Venice"

%
Jag somnade läsa en tråkig bok, och jag drömde att jag läste på,så jag vaknade upp från ren tristess.
		-- William Shakespeare, "The Merchant of Venice"

%
Jag har aldrig låta min skolgång störa med min utbildning.
		-- Mark Twain

%
Jag måste ha en ofantlig mängd sinnes; det tar mig så mycket som envecka ibland för att göra upp.
		-- Mark Twain, "The Innocents Abroad"

%
Jag tror vördnads att tillverkaren som gjorde oss alla gör allt i NewEngland, men vädret. Jag vet inte vem som gör det, men jag tror att det måste vararåa lärlingar i väder kontorister fabrik som experiment och lära sig hur, iNew England, för kost och kläder, och sedan främjas för att göra väder förländer som kräver en bra artikel, och kommer att ta deras sed på annat hållom de inte får det.
		-- Mark Twain

%
Jag tror att vi är i råttornas Alley där de döda män förlorat sina ben.
		-- T.S. Eliot

%
Jag var glada att kunna svara snabbt, och jag gjorde. Jag sa att jag inte visste.
		-- Mark Twain

%
Jag kommer att hedra julen i mitt hjärta, och försöker hålla det hela året. jagkommer att leva i det förflutna, nutid och framtid. Andar allaTre skall sträva inom mig. Jag kommer inte att stänga ute de lärdomar som delära. Åh, säg att jag kan svamp bort skriften på denna sten!
		-- Charles Dickens

%
"Jag undrar", sade han till sig själv, "vad som finns i en bok medan den är stängd. Åh, jagvet att det är fullt av bokstäver tryckta på papper, men i alla fall, något måstehända, eftersom så fort jag öppnar det, det finns en hel berättelse med människorJag vet inte ännu och alla typer av äventyr och strider. "
		-- Bastian B. Bux

%
Jag ska bränna mina böcker.
		-- Christopher Marlowe

%
Jag har touch'd den högsta punkten av hela mitt storhet;Och från att full meridianen min äraJag skynda nu till min inställning. Jag skall falla,Som en ljus utandning på kvällenOch ingen människa kan se mig mer.
		-- Shakespeare

%
Om fler av oss värderas mat och jubel och sång ovan hamstrade guld, skulle detvara en desto bättre världen.
		-- J.R.R. Tolkien

%
Om man inte kan njuta av att läsa en bok om och om igen, det är ingen idéläsa det alls.
		-- Oscar Wilde

%
Om två människor älskar varandra, kan det inte finnas någon lyckligt slut för det.
		-- Ernest Hemingway

%
Om du som alla våra lagar början till slut, skulle det inte finnas något slut.
		-- Mark Twain

%
Om du plockar upp en svältande hund och gör honom välmående, kommer han inte bita dig.Detta är den huvudsakliga skillnaden mellan en hund och en man.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Om du berättar sanningen du inte behöver komma ihåg något.
		-- Mark Twain

%
I ett museum i Havanna, det finns två skallar av Christopher Columbus,"En när han var en pojke och en när han var en människa."
		-- Mark Twain

%
I Indien, "kallt väder" är bara en vanlig fras och har kommit inanvända genom nödvändigheten av att ha något sätt att skilja mellan vädersom kommer att smälta en mässingsdörrvredet och väder som endast kommer att göra det mosig.
		-- Mark Twain

%
I Marseille gör de halva toalettvål vi konsumerar i Amerika, menMarseljäsen har bara en vag teoretisk uppfattning om dess användning, som dehar erhållits från böcker av resor.
		-- Mark Twain

%
För det första, gjorde Gud idioter; Detta var för att öva; sedan gjorde hanskolstyrelser.
		-- Mark Twain

%
I handlingen, folk kom till landet; landet älskade dem; de arbetade ochkämpade och hade massor av barn. Det var en fransman som talade roligoch en gröngöling från England som var en fancy-pants men när det kom tillkritan han var allt mod. Dessa romaner skulle göra dig kväljningar.roman.
		-- Canadian novelist Robertson Davies, on the generic Canadian

%
Inom loppet av ett hundra sjuttiosex år Mississippi harförkortas sig två hundra fyrtiotvå miles. Därför ... i GamlaSilur Period Mississippifloden var uppåt en miljon trehundratusen miles lång ... sjuhundra fyrtiotvå år från nuMississippi blir bara en mil och tre fjärdedelar lång. ... Det finnsnågot fascinerande om vetenskap. Man får sådana hälso avkastninggissningar ur en sådan obetydlig investering på faktum.
		-- Mark Twain

%
Under våren har jag räknade 136 olika typer av väder inuti24 timmar.
		-- Mark Twain, on New England weather

%
Det har länge varit ett axiom av min som de små saker är oändligtdet viktigaste.
		-- Sir Arthur Conan Doyle, "A Case of Identity"

%
Det är en klok far som känner sitt eget barn.
		-- William Shakespeare, "The Merchant of Venice"

%
Det är genom turen att Gud att i det här landet, har vi tre fördelar:yttrandefrihet, tankefrihet, och visdom aldrig att använda antingen.
		-- Mark Twain

%
Det är lätt att hitta fel, om man har det disposition. Det var en gång en mansom att inte kunna hitta någon annan fel med sin kol, klagade över attdet fanns alltför många förhistoriska paddor i det.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Det är ofta fallet att man som inte kan ljuga tror att han är den bästadomare en.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Det är rätt att han också skulle ha sin lilla krönika, sina minnen,hans skäl, och kunna känna igen det goda i det dåliga, dåligt ivärst, och så växer försiktigt gammal alla ned oföränderliga dagar och dö endag som alla andra dagar, bara kortare.
		-- Samuel Beckett, "Malone Dies"

%
Det tar oftast mer än tre veckor att förbereda ett bra improviserat tal.
		-- Mark Twain

%
Det var inte det bästa som vi alla bör tänka lika; det är meningsskiljaktighetersom gör hästkapplöpningar.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Dess namn är den allmänna opinionen. Den hålls i vördnad. Det avgör allt.Vissa tycker att det är Guds röst.
		-- Mark Twain

%
Vänlighet är ett språk som döva kan höra och blinda kan läsa.
		-- Mark Twain

%
Kiss me, Kate, kommer vi att vara gifta o söndag.
		-- William Shakespeare, "The Taming of the Shrew"

%
Låg på, MacDuff och curs'd vara den som först ropar, "Hold, nog!".
		-- Shakespeare

%
Låt honom välja ut mina filer, hans projekt att åstadkomma.
		-- Shakespeare, "Coriolanus"

%
Låt mig ta dig en knapp-hål lägre.
		-- William Shakespeare, "Love's Labour's Lost"

%
Låt oss sträva efter att leva på att när vi kommer att dö även begravnings blirförlåt.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Som en dyr sportbil, finjusteras och välbyggd, Portia var snygg,välväxt och vacker, hennes röda overall gjutning hennes kropp, som var så varmsom seatcovers i juli håret så mörk som nya däck, hennes ögon blinka somljusa navkapslar, och hennes läppar som daggiga som pärlorna av färsk regn på huven;Hon var en kvinna som drivs - drivs av en enda accelerator - och hon behövde enman, en man som inte skulle flytta från sina vyer, en man att styra henne längsrätt väg: en man som Alf Romeo.Håret bollen blockerar avloppet i duschen påminde Laura hon skulle aldrigse hennes lilla hund Pritzi igen.Det kunde ha varit en organiskt baserad störning i hjärnan - kanske entumör eller en metabolisk brist - men efter en grundlig neurologisk undersökning detbestämdes att Byron var helt enkelt en idiot.Vinnare i den 7: e årliga Bulwer-Lytton Bad Writing Contest. Tävlingen äruppkallad efter författaren till de odödliga rader: "Det var en mörk och stormignatt. "Syftet med tävlingen är att skriva den första meningen i detsämsta möjliga roman.
		-- Jeff Jahnke, runner-up

%
Herre, vad bedrar dessa dödligar!
		-- William Shakespeare, "A Midsummer-Night's Dream"

%
Människan är det enda djur som rodnar - eller behöver.
		-- Mark Twain

%
Många författare verkar tro att han är aldrig djup utom när han inte kanförstå sin egen mening.
		-- George D. Prentice

%
Många rasande psykiatriker anstiftan en trött slaktare. Slaktaren ärtrötta och trött eftersom han har styckat kött och stek och lamm i timmar ochveckor. Han önskar inte att sjunga om något med raving psykiatriker,men han sjunger om sin gingivectomist, han drömmer om en enda cosmologist,han tycker om sin hund. Hunden heter Herbert.
		-- Racter, "The Policeman's Beard is Half-Constructed"

%
Många sidor gör en tjock bok, med undantag för fick biblar som är på mycketmycket tunt papper.
		-- Racter, "The Policeman's Beard is Half-Constructed"

%
Många sidor gör en tjock bok.
		-- Racter, "The Policeman's Beard is Half-Constructed"

%
Sinne! Jag menar inte att säga att jag vet, min egen kunskap, vad som finnssärskilt död om en dörr-spik. Jag kan ha lutande själv,att betrakta en kista-spik som deadest bit beslag i handeln.Men visdom våra förfäder är i liknelse; och mina ohelig händerfår inte störa den, eller landets gjort för. Du kommer därför tillåtamig att upprepa, med eftertryck, att Marley var lika död som en dörr spik.
		-- Charles Dickens, "A Christmas Carol"

%
Måste jag hålla ett ljus till mina shames?
		-- William Shakespeare, "The Merchant of Venice"

%
Mina kära människor.Min kära Bagginses och Boffins, och min kära Tooks och Brandybucks,och Grubbs, och Chubbs, och Burrowses, och Hornblowers och Bolgers,Bracegirdles, Goodbodies, Brockhouses och Proudfoots. Också min godaSack Bagginses att jag välkommen tillbaka äntligen Bag End. Idag är min111:e födelsedag: Jag är eleventy-en dag "!
		-- J. R. R. Tolkien

%
Min enda kärlek sprungen ur min enda hat!För tidigt sett okända och kända för sent!
		-- William Shakespeare, "Romeo and Juliet"

%
skrattar aldrig på levande drakar.
		-- Bilbo Baggins [J.R.R. Tolkien, "The Hobbit"]

%
Ingen grupp av personal möter utom att konspirera mot den breda allmänheten.
		-- Mark Twain

%
Inga levande organism kan fortsätta under lång tid att existera förnuftigt under förhållanden medabsolut verklighet; även lärkor och katydids är tänkt, av vissa, att drömma.Hill House, inte frisk, stod sig mot sina kullar, hålla mörkretinom; det hade stått så i åttio år och kan stå för åttio mer.Inom väggar fortsatt upprätt, tegel möttes snyggt, golv var fast, ochdörrar förnuftigt stängdes; tystnad låg stadigt mot trä och stenav Hill House, och vad gick det, gick ensam.
		-- Shirley Jackson, "The Haunting of Hill House"

%
Inget våld, mina herrar - inget våld, jag ber dig! Tänk på möbler!
		-- Sherlock Holmes

%
Buller bevisar ingenting. Ofta en höna som bara har lagt ett ägg kacklarsom om hon lade en asteroid.
		-- Mark Twain

%
"Inte Hercules kunde ha knock'd ut sina hjärnor, för han hade ingen."
		-- Shakespeare

%
Ingenting så behöver reformeras som andras vanor.
		-- Mark Twain

%
Ingenting så behöver reformeras som andras vanor.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
O, det är utmärktAtt ha en jätte styrka; men det är tyranniskFör att använda den som en jätte.
		-- Shakespeare, "Measure for Measure", II, 2

%
12 oktober Discovery.Det var underbart att hitta Amerika, men det skulle ha varit mer underbart att missaDet.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Oktober.Detta är en av de säregna farliga månader att spekulera i aktier i.De andra är juli, januari, September, April, November, maj, mars, juni,December, augusti och februari.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
O, vad en tilltrasslad webb vi väver, när först vi övar att bedra.
		-- Sir Walter Scott, "Marmion"

%
En av de mest slående skillnaderna mellan en katt och en lögn är att en katt harbara nio liv.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Patch sorger med ordspråk.
		-- William Shakespeare, "Much Ado About Nothing"

%
Farlig för oss alla är de enheter av en konst djupare än vi självabesitter.
		-- Gandalf the Grey [J.R.R. Tolkien, "Lord of the Rings"]

%
Personer som försöker att hitta ett motiv i denna berättelse kommer att åtalas;personer som försöker att hitta en moralisk i den kommer att förvisas; personer som försökeratt hitta en tomt i det kommer att skjutas. Genom beslut av författaren
		-- Mark Twain, "The Adventures of Huckleberry Finn"

%
fråga = (till)? vara:! vara;
		-- Wm. Shakespeare

%
Reader Anta att du var en idiot. Och antar att du var en medlem avKongress. Men jag upprepar mig.
		-- Mark Twain

%
Rebellion låg i hans väg, och han fann det.
		-- William Shakespeare, "Henry IV"

%
Anmärkning av Dr Baldwins om uppkomlingar: Vi bryr oss inte att äta svamparsom tror att de är tryffel.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Repliker är något vi tänker på tjugofyra timmar för sent.
		-- Mark Twain

%
ROMEO: Mod, man; ont kan inte vara mycket.Mercutio: Nej, 'tis inte så djupt som en brunn, eller så bredsom en kyrkdörren; men 'tis nog, "twill tjäna.
		-- Mark Twain

%
Att se till att död, en nödvändig ände,Kommer när det kommer.
		-- William Shakespeare, "Julius Caesar"

%
Hon är raffinerade. Hon är inte oraffinerad. Hon håller en papegoja.
		-- Mark Twain

%
Sheriff Chameleotoptor suckade med en air av trötta sorg, och sedanvände sig till Doppelgutt och sade "Senator måste verkligen ha varit på enBender här gången - han lämnade en fest i Cleveland, Ohio, på 11:30 sistanatten, och de hittade hans bil i morse i skorstenen av en brittiskhangarfartyg i Formosa Straits. "dålig fiction tävling.
		-- Grand Panjandrum's Special Award, 1985 Bulwer-Lytton

%
Små saker gör bas män stolt.
		-- William Shakespeare, "Henry VI"

%
Så gick hon ut i trädgården för att skära en kål blad för att göra en äppelpaj;och samtidigt en stor björninna, som kommer upp på gatan dyker huvudetin i butiken. "Vad! Ingen tvål?" Han dog, och hon mycket oförsiktigtgift barberaren; och det fanns närvarande Picninnies och GrandSMÅPÅVE själv, med den lilla runda knappen längst upp, och allaföll till att spela spelet fångst som fångst kan, tills krut sprangut på hälarna på sina stövlar.
		-- Samuel Foote

%
Så så är bra, mycket bra, mycket bra bra:och ändå är det inte; det är men så så.
		-- William Shakespeare, "As You Like It"

%
Tvål och utbildning är inte lika plötsligt som en massaker, men de är merdödligt i det långa loppet.
		-- Mark Twain

%
Något är ruttet i staten Danmark.
		-- Shakespeare

%
Ibland undrar jag om jag i min högra sinne. Då den passerar ut och jag ärlika intelligent som någonsin.
		-- Samuel Beckett, "Endgame"

%
"Säg, du vast och anrika huvudet," muttrade Ahab ", som, ävenungarnished med ett skägg, men här och där lookest hoary med mossa; tala,mäktig huvud, och berätta hemligheten sak som är i dig. Av alla dykare,du har dykt djupare. Att huvudet på vilken den övre sön glimmar nu harflyttade mitt världens grundvalar. Där oregistrerade namn och flottor rostar,och outsägligt hopp och ankare ruttna; där i hennes mord hålla denna fregattJorden ballast med ben miljoner av drunknade; där, i den fruktansvärdavatten-land, det var din mest kända hem. Du har varit där klocka ellerdykare gick aldrig; har sovit med många seglare sida, där sömnlösa mödrarskulle ge sina liv för att fastställa dem. Thou saw'st de låsta älskande närhoppar från deras brinnande fartyg; hjärta till hjärta de sjönk under triumferarvåg; trogna varandra, när himlen verkade falska dem. Thou saw'st denmördade mate när kastas av pirater från midnatt däck; timmar han föllin i den djupare midnatt av OMÄTTLIG gap; och hans mördare fortfarande segladepå oskadda - medan snabba blixtar ryste grann fartyget som skullehar burit en rättfärdig man att utsträckt, längtande armar. O huvud! thou harsett tillräckligt för att dela planeterna och göra en otrogen Abrahams, och inte enstavelse är ditt! "
		-- H. Melville, "Moby Dick"

%
Stadig rörelse är viktigare än hastighet, mycket av tiden. Så längeeftersom det finns en regelbunden progression av stimuli för att få din mentala krokarin i, det finns utrymme för rörelse i sidled. När detta börjar, är dess hastigheten fråga om bedömning.
		-- Corwin, Prince of Amber

%
Sluta! Det var först en omgång Blindman bock. Naturligtvis fanns.Och jag inte mer tror Topper var verkligen blinda än jag tror att han hade ögoni sina stövlar. Min uppfattning är att det var en klar sak mellan honom ochScrooges systerson, och att spöken av julklapp visste det. Dehur han gick efter det knubbig syster i spets Tucker, var en skandalpå godtrogenhet av den mänskliga naturen.
		-- Corwin, Prince of Amber

%
Misstanke hemsöker alltid de skyldiga sinnet.
		-- Wm. Shakespeare

%
Swerve mig? Vägen till min fasta syfte läggs med järnskenor,varpå min själ räfflad att köra. Över unsounded raviner, genomde plundrade hjärtan berg, under enter "sängar, ofelbart jag rusa!
		-- Captain Ahab, "Moby Dick"

%
Talare finns inga bra doers.
		-- William Shakespeare, "Henry VI"

%
Tala sanning eller trumf - men få tricket.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Fresta inte ett desperat man.
		-- William Shakespeare, "Romeo and Juliet"

%
Missbruket av storheten är när det disjoins ånger från makten.
		-- William Shakespeare, "Julius Caesar"

%
Viken-träd i vårt land är alla wither'dOch meteorer skrämsel de fasta stjärnorna på himmelen;Den bleka månen ser blodiga på jordenOch lean-look'd profeter viska rädda förändring.Dessa tecken förfraktion död eller hösten kungar.
		-- Wm. Shakespeare, "Richard II"

%
Den större delen av tapperhet är diskretion.
		-- William Shakespeare, "Henry IV"

%
Den iskall skrik dela den varma sommarnatten i två, den förstahälften är före skrik när det var ganska ljumma och lugn ochtrevlig, andra hälften fortfarande ljumma och ganska trevlig för dem somhade inte hört skrik alls, men inte lugn eller ljumma eller till och med mycket trevligför dem som hörde skrik, diskontera den lilla tidunder själva skrika sig när dina öron kanske har hört detmen din hjärna inte reagera ännu så att du vet.
		-- Winning sentence, 1986 Bulwer-Lytton bad fiction contest.

%
Den Bulwer-Lytton fiktion tävling hålls någonsin år på San Jose StateUniv. av professor Scott Rice. Den hålls till minne av Edward GeorgeEarle Bulwer-Lytton (1803-1873), en ganska produktiv och populär (i hanstid) författaren. Han är mest känd idag för att ha skrivit "The LastDagar av Pompeji. "När Snobben börjar skriva sin roman från toppen av sin hundkoja,början "Det var en mörk och stormig natt ..." han lånar från LordBulwer-Lytton. Detta var den linje som öppnade sin roman, "Paul Clifford,"skriven i 1830. Den fullständiga linjen avslöjar varför det är så illa:Det var en mörk och stormig natt; regnet föll i strömmar - utomvid tillfälliga intervaller, när den kontrollerades av en våldsam pust avvind som svepte upp gatorna (för det är i London som vår scenligger), skramlande längs hustaken, och häftigt röra om knapphändigaflamma av lamporna som kämpade mot mörkret.
		-- Winning sentence, 1986 Bulwer-Lytton bad fiction contest.

%
Kamelen dog helt plötsligt på den andra dagen, och Selena frettedtrumpet och putsning henne redan oklanderlig naglar - inte för förstagången sedan resan begain - funderade snidely om detta skulle lösa uppi en vinjett av mindre besvär som alla andra helgdagar tillbringademed basilika.
		-- Winning sentence, 1983 Bulwer-Lytton bad fiction contest.

%
Nedräkningen hade stannat vid "T" minus 69 sekunder när Desiree, den förstakvinnlig apa att gå upp i rymden, blinkade åt mig slugt och tjurade hennes tjocka,gummi läppar otvetydigt - den första av många sådana framsteg under detskulle visa sig vara den längsta och mest minnesvärda, rymdfärden minkarriär.
		-- Winning sentence, 1985 Bulwer-Lytton bad fiction contest.

%
Djävulen kan citera Skriften för hans ändamål.
		-- William Shakespeare, "The Merchant of Venice"

%
Skillnaden mellan ett mirakel och en Faktum är exakt skillnadenmellan en sjöjungfru och en tätning.
		-- Mark Twain

%
Skillnaden mellan det rätta ordet och den nästan rätt ord är denskillnaden mellan blixt och blixten bug.
		-- Mark Twain

%
Mode bär mer kläder än mannen.
		-- William Shakespeare, "Much Ado About Nothing"

%
Det första vi gör, låt oss döda alla advokater.
		-- Wm. Shakespeare, "Henry VI", Part IV

%
Den heliga passion Vänskap är så söt och stadig och lojal ochvaraktig natur att det kommer att pågå igenom en hel livstid, om inte begärt attlåna pengar.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Den mänskliga rasen har ett riktigt effektivt vapen, och det är skratt.
		-- Mark Twain

%
Den mänskliga rasen är en ras av ynkryggar, och jag är inte bara marscherar i detprocession men bär en banderoll.
		-- Mark Twain

%
Det sista man vet att konstruera ett verk är vad man ska sätta först.
		-- Blaise Pascal

%
Least Lyhörd litteraturkritikerDen viktigaste kritiker i vårt område av studien är Lord Halifax. enmest individuella domare poesi, han en gång bjöd Alexander Pope runt tillge en offentlig läsning av hans senaste dikt.Pope, ledande poet av hans dag, blev mycket förvånad när LordHalifax stoppade honom fyra eller fem gånger och sa, "Jag ber om ursäkt, Mr.Pope, men det finns något i den passage som inte riktigt tillfredsställa mig. "Pope gjordes mållös, eftersom detta fina kritiker föreslog betydandeoch okloka emendations till hans senaste mästerverk. "Var så god och markeraplatsen och överväga på din fritid. Jag är säker på att du kan ge det en bättresväng."Efter läsningen, en god vän till Lord Halifax, en viss Dr.Garth tog bedövade påven åt sidan. "Det finns inget behov av att röralinjer ", sade han." Allt du behöver göra är att lämna dem precis som de är, uppmanaLord Halifax två eller tre månader därmed, tacka honom för hans vänliga observationpå dessa avsnitt, och sedan läsa dem till honom som ändras. Jag har känt honommycket längre än du har, och kommer att vara ansvarig för händelsen. "Påven tog hans råd, uppmanade Lord Halifax och läste diktenprecis som det var innan. Hans unika kritiska förmåga hade förlorat något avderas kant. "Ay", kommenterade han, "nu är de helt rätt. Ingenting kanbli bättre."
		-- Stephen Pile, "The Book of Heroic Failures"

%
Den minst framgångsrika CollectorBetsy Baker spelade en central roll i historien att samla in. Honanvändes som en tjänare i huset av John Warburton (1682-1759) som hadesamlat en fin samling av 58 första upplagan pjäser, däribland de flesta avverk av Shakespeare.En dag Warburton återvände hem för att hitta 55 av dem förkolnade bortomläsbarhet. Betsy hade antingen brände dem eller använt dem som en plätt bottnar. Deåterstående tre folios är nu i British Museum.Den enda jämförbara litterära figur var maid som i 1835 brannmanuskriptet till den första volymen av Thomas Carlyle "The Hisory avFranska revolutionen ", tänkte att det var returpapper.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Den vackra flickebarn Kaa var obarmhärtigt kedjad till den grymma postenkrigaren chefredaktör Beast, med sin barbar stam nu stapla ved påhennes nubile fötter, när den starka tydlig röst poetiska och heroiskaHandsomas röt, 'snärta din Bic, skarpa att chick, och du kommer att känna minstål genom din sista måltid! "
		-- Winning sentence, 1984 Bulwer-Lytton bad fiction contest.

%
Galningen, älskaren och poeten,Är fantasi alla kompakta ...
		-- Wm. Shakespeare, "A Midsummer Night's Dream"

%
Mannen som syftar till att göra en katt med svansen lär sig något somkommer alltid att vara användbar och som aldrig kommer att växa svag eller tveksam.
		-- Mark Twain

%
Den nakna sanningen om det är, jag har ingen skjorta.
		-- William Shakespeare, "Love's Labour's Lost"

%
"... Namnet på låten heter" Haddocks 'Eyes'! ""Åh, det är namnet på låten, är det?" Alice sa, försökerkänner dig intresserad."Nej, du förstår inte" riddaren sade, ser liteförargad. "Det är vad namnet heter. Namnet verkligen är," The AgedMedelålders man. ""Då jag borde ha sagt" Det är vad låten heter "?"Alice korrigerade sig."Nej, du borde inte: det är en helt annan sak Låten ärkallade ways and means ", men det är bara vad det kallas du vet"!"Nå, vad är låten då?" sade Alice, som var av dennatid förvirrade helt."Jag var på väg till det", sade riddaren. "Låten är verkligen"A-sitter på en Gate" och låten är min egen uppfinning ".
		-- Lewis Carroll, "Through the Looking Glass"

%
Noterna blatted mot himlen när de steg över Kanada gäss, befjädradegump mooning dagen, simhud bihang frenetiskt trampa oseddacyklar i sitt sökande efter näring, som drivs av grym naturens maxim,"Ya vill äta, ya gotta arbete," och till sist jag visste Pittsburgh.
		-- Winning sentence, 1987 Bulwer-Lytton bad fiction contest.

%
De enda människor för mig är galna som - de som är galna att leva,galna att prata, galna som ska sparas, önskar allt på samma gång,de som aldrig gäspa eller säga en vanlig sak, men bränna, bränna, brännasom fantastiska gula romerska ljus.
		-- Jack Kerouac, "On the Road"

%
Det enda sättet att hålla din hälsa är att äta vad du inte vill, dricka vaddu inte gillar, och gör vad du inte vill.
		-- Mark Twain

%
Prästens grå nimbus i en nisch där han klädd diskret.Jag kommer inte att sova här i kväll. Hem också jag kan inte gå.En röst, sötad och ihållande, ropade på honom från havet.Vrida kurvan han vinkade med handen. En elegant brunt huvud, en säl, långtut på vattnet, runda. Inkräktare.
		-- James Joyce, "Ulysses"

%
Allmänheten är bara en multiplicerad "mig."
		-- Mark Twain

%
Den mognaste frukten faller först.
		-- William Shakespeare, "Richard II"

%
Hemligheten källa för humor är inte glädje men sorg; det finns ingen humor i himlen.
		-- Mark Twain

%
Den minsta mask blir att trampas på.
		-- William Shakespeare, "Henry VI"

%
Det säkraste skyddet mot frestelsen är feghet.
		-- Mark Twain

%
Den sanna södra vattenmelon är en välsignelse varandra, och inte nämnas medvanligare saker. Det är chef för världens lyx, kung av Guds nådöver alla frukterna av jorden. När man har ätit det, vet vad hanänglar äter. Det var inte en sydlig vattenmelon att Eva tog; Vi vet det eftersomhon omvände.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Själva bläck med vilken all historia skrivs är bara vätska fördomar.
		-- Mark Twain

%
Det finns fler saker i himmel och jord,Horatio, än är drömt om i din filosofi.
		-- Wm. Shakespeare, "Hamlet"

%
Det finns tre ofelbara sätt att talande en författare, och tre bildar enstigande skala av komplimang: en, för att tala om för honom att du har läst en av hans böcker; 2,att berätta för honom att du har läst alla hans böcker; 3, för att be honom att låta dig läsamanuskriptet till sin kommande bok. Nr 1 medger dig till sin respekt; No. 2medger du att hans beundran; Nr 3 bär dig klar i hans hjärta.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Det finns en stor upptäckt fortfarande göras i litteratur: attbetala litterära män av den kvantitet som de inte skriver.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Det finns alltid en sak att komma ihåg: författare alltid säljer någon ut.
		-- Joan Didion, "Slouching Towards Bethlehem"

%
Det finns en gammal tid toast som är gyllene för sin skönhet."När du uppför kullen välstånd kan du inte träffa en vän."
		-- Mark Twain

%
Det finns inget tecken, oavsett hur bra och bra, men det kan förstöras avförlöjliga, oavsett hur dålig och dum. Observera röven, till exempel: hanstecken om perfekt, är han de ädlaste andan bland alla humblerdjur, men se vad förlöjligande har fört honom till. I stället för känslakompletterat när vi kallas en åsna, vi kvar i tvivel.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Det finns ingen distinkt indian kriminell klass utom kongressen.
		-- Mark Twain

%
Det finns ingen jakt som jakt på mannen, och de som har jagatbeväpnade män tillräckligt länge och gillade det, aldrig ta hand om något annat därefter.
		-- Ernest Hemingway

%
Det finns små val i ruttna äpplen.
		-- William Shakespeare, "The Taming of the Shrew"

%
De har varit på en stor fest språk, och stulna resterna.
		-- William Shakespeare, "Love's Labour's Lost"

%
De stava det "da Vinci" och uttalas "da Vinchy". utlänningaralltid stava bättre än de uttala.
		-- Mark Twain

%
Saker tidigare prövning och nu med mig förbi vård.
		-- William Shakespeare, "Richard II"

%
Detta är den första ålders som är ägnat mycket uppmärksamhet åt framtiden, vilket är enlite ironiskt eftersom vi inte kan ha en.
		-- Arthur Clarke

%
Denna natt methinks är bara dagsljus sjuka.
		-- William Shakespeare, "The Merchant of Venice"

%
Detta var den mest unkindest skära av alla.
		-- William Shakespeare, "Julius Caesar"

%
Att vara eller inte vara.Att göra är att vara.Att vara är att göra.Gör att göra att göra.
		-- Sinatra

%
För mycket är lagom.
		-- Mark Twain, on whiskey

%
Utbildning är allt. Peach var en gång en bittermandel; blomkål äringenting men kål med en högskoleutbildning.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Sanningen är det mest värdefulla vi har - så låt oss hushålla det.
		-- Mark Twain

%
Såvida timmar var koppar säck, och minuter kapuner, och klockar tungornaav bawds, och rattar tecken på hoppande hus, och välsignade solen självett rättvist, varm wench i flamma-färgad taft, ser jag ingen anledning till varför du skallvara så överflödigt att kräva tid på dagen. Jag slöseri med tid och nu dothtid avfall mig.
		-- William Shakespeare

%
Wagners musik är bättre än det låter.
		-- Mark Twain

%
Vatten, tas med måtta kan inte skada någon.
		-- Mark Twain

%
Vi vet allt om vanor myran, vi vet allt om vanorbee, men vi vet ingenting alls om vanor ostron. Det verkarnästan säker på att vi har valt fel tidpunkt för att studeraostron.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Vi bör vara noga med att ta sig ur en upplevelse bara visdom som äri det - och stanna där, så att vi som katten som sätter sig på en varmspis-lock. Hon kommer aldrig att sitta på en het spis-locket igen - och attär väl; men också att hon aldrig kommer att sitta på en kall längre.
		-- Mark Twain

%
Vi var unga och vår lycka bländas oss med sin styrka. Men det fannsockså ett fruktansvärt svek som låg inom mig som en Merle Haggard låten på enFransk restaurang. [...]Jag kunde inte berätta flickan om kvinnan i tollway, hennes mjölkvit BMW och hennes Jordache leende. Det hade varit en kamp. Jag hade stansade hennepojkvän, som kämpade mot mekanisk tjur. Alla sa till honom: "Du ridatjur, senor. Du behöver inte bekämpa den. "Men han var mager och hård som en dåligrib-ögat och han kämpade tjuren. Och då han kämpade mig. Och när vi avslutatDet fanns inga vinnare, bara män gör vad män måste göra. [...]"Stanna bilen", sade flickan.Det var en blick av fruktansvärd sorg i ögonen. Hon kände tillkvinna tollway. Jag visste inte hur. Jag började tala, men hon höjde ettarm och talade med en lugn och frid som jag aldrig kommer att glömma."Jag ber inte om vem är tollway belle", sade hon, "tollwayBelle för dig. "Nästa morgon våra ungdomar var ett minne, och vår lycka var en lögn.Livet är som en dålig margarita med bra tequila, jag tänkte som jag hällde whiskypå min granola och inför en ny dag.konkurrens
		-- Peter Applebome, International Imitation Hemingway

%
Hur som helst, jag läser detta James Bond bok, och genast insåg jagdet som de flesta böcker, hade det alltför många ord. Handlingen var densamma somalla James Bond böcker har: En ond person försöker att spränga världen, menJames Bond dödar honom och hans hantlangare och gör kärlek till flera attraktivakvinnor. Där det är det: 24 ord. Men killen som skrev boken tog* tusentals * ord att säga det.Eller tänk "Bröderna Karamazov", den berömda ryska alkoholFjodor Dostojevskij. Det handlar om dessa två bröder som dödar sin far.Eller kanske bara en av dem dödar fadern. Det är omöjligt att säga eftersomvad de oftast gör är att prata för nästan tusen sidor. Om alla ryssar pratalika mycket som Karamazovs gjorde, jag kan inte se hur de funnit tid att bli enstormakt.Man säger att Dostojevskij skrev "Bröderna Karamazov" för att höjaFrågan om huruvida det finns en Gud. Varför kom han inte bara rättut och säga: "Finns det en Gud Det slår säkert heck av mig?".Andra kända verk kunde lätt har sammanfattats i ett par ord:* "Moby Dick" - Bråka inte runt med stora valar eftersom de symboliserar  natur och kommer att döda dig.* "Två städer" - fransmän är galna.
		-- Dave Barry

%
Hur bra är en obscenitet rättegången förutom att popularisera litteratur?
		-- Nero Wolfe, "The League of Frightened Men"

%
Vad jag berätta tre gånger är sant.
		-- Lewis Carroll

%
Vad ingen make till en författare någonsin kan förstå är att en författare arbetarnär han stirrar ut genom fönstret.
		-- Lewis Carroll

%
När arg, räkna fyra; när mycket arg, svär.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
När jag tänker på antalet obehag människor som jag känner som har gåtttill en bättre värld, jag flyttade till leva ett annat liv.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
När jag var yngre, jag kunde komma ihåg något, om det hade hänteller inte; men mina fakulteter ruttnande nu och jag ska snart vara så jagkan inte komma ihåg något, men de saker som aldrig hänt. Det är tråkigt attgå sönder så här men vi alla måste göra det.
		-- Mark Twain

%
När du är osäker, tala sanning.
		-- Mark Twain

%
När en bränner sina broar, vad en mycket trevlig brand det gör.
		-- Dylan Thomas

%
När du är på väg att dö, är en wombat bättre än inget företag alls.
		-- Roger Zelazny, "Doorways in the Sand"

%
Närhelst litterära tyska dyk i en mening, är att den sistadu kommer att se av honom tills han dyker upp på den andra sidan av hansAtlanten med sin verb i munnen.
		-- Mark Twain "A Connecticut Yankee in King Arthur's Court"

%
När du upptäcker att du är på sidan av majoriteten, är det dagsatt reformera.
		-- Mark Twain

%
Den som har levt tillräckligt länge för att ta reda på vad livet är, vet hur djupt en skuldtacksamhet vi är skyldiga till Adam, den första stora välgörare vår ras. hanförde död i världen.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Varför är det så att vi glädjas åt en förlossning och sörjer vid en begravning? Det beror på att viär inte den berörda personen.
		-- Mark Twain, "Pudd'nhead Wilson's Calendar"

%
Arbetet består av vad en kropp är skyldig att göra.Spela består av vad en kropp inte är skyldig att göra.
		-- Mark Twain

%
Rynkor bör endast ange var leenden har varit.
		-- Mark Twain

%
Att skriva är lätt; allt du behöver göra är att sitta stirrar på tomt pappersark tillsdroppar blod formulär på din panna.
		-- Gene Fowler

%
Skrift vänder sina värsta stunder i pengar.
		-- J.P. Donleavy

%
"Du har varit i Afghanistan, jag uppfattar."
		-- Sir Arthur Conan Doyle, "A Study in Scarlet"

%
"Ni har hört mig tala om professor Moriarty?""Den berömda vetenskapliga brottsling, lika känd bland skurkar som -""Mina rodnar, Watson," Holmes mumlade, i en avvärjande röst."Jag var på väg att säga" som han är okänd för allmänheten. "
		-- A. Conan Doyle, "The Valley of Fear"

%
Du kanske mina härligheter och mitt tillstånd avyttra,Men inte mina sorger; fortfarande är jag kung av dem.
		-- William Shakespeare, "Richard II"

%
Ni nämnde ditt namn som om jag skulle känna igen det, men utöver detuppenbara fakta som du är en kandidat, en advokat, en frimurare, ochen astmatiker, jag vet ingenting alls om dig.
		-- Sherlock Holmes, "The Norwood Builder"

%
Du behöver aldrig ändra något du fick upp mitt i nattenatt skriva.
		-- Saul Bellow

%
Du ser, jag anser att en människas hjärna ursprungligen är som en liten tomtvinden, och man måste fylla på med sådana möbler som du väljer. En dåretar in all bråte av varje slag han kommer över, så att kunskapensom kan vara till nytta för honom blir trångt ut, eller i bästa fall är konfys meden hel del andra saker, så att han har svårt att lägga sina händer på det.Nu skicklig arbetare är mycket försiktig verkligen vad han tar i sinbrain-vinden. Han kommer att ha något annat än de verktyg som kan hjälpa honom att görahans arbete, men av dessa har han ett stort sortiment, och alla i den mest perfektabeställa. Det är ett misstag att tro att det lilla rummet har elastiska väggar ochkan tänja i någon utsträckning. Beroende på den det kommer en tid då för varjeFörutom kunskap du glömmer något som du visste innan. Den är avstörsta vikt, därför att inte ha onödiga fakta att inverkade användbara sådana.
		-- Sir Arthur Conan Doyle, "A Study in Scarlet"

%
Du beträder mitt tålamod.
		-- William Shakespeare, "Henry IV"

%
Ni minns, Watson, hur fruktansvärda verksamheten iAbernetty familj först kom till min kännedom av djupet sompersilja hade sjunkit i smöret på en varm dag.
		-- Sherlock Holmes

%
Ditt manus är både bra och originell, men den del som är bra är inteoriginal och den del som är original är inte bra.
		-- Samuel Johnson

%
Zounds! Jag var aldrig så bethumped med ordeftersom jag först ringde min brors pappa pappa.
		-- William Shakespeare, "Kind John"

%
Sinnet är sin egen plats, och i sigKan göra en Him'len Hell, ett helvete av Him'len.
		-- John Milton

%
"Jag förstår att detta är din första döda klient" Sabian sade. Deabsurda i uttalandet jag vill skratta men de inte kalla migUttryckslöst Allie och lögn.
		-- Pat Cadigan, "Mindplayers"

%
En bårhuset är ett bårhus är ett bårhus. De kan måla väggarna med aggressivtglada grundfärger och splashy snygg grafik, men det är fortfarande en anläggningplats för de döda tills de kan skiljas ut till banker organ. Inte för att jagskulle ha omhändertagna normalt men min synvinkel var skev. den obevekligaPleasence av rummet jag satt i verkade bara groteskt.
		-- Pat Cadigan, "Mindplayers"

%
"Vad är det här Trix? Tant! Trix? Dig? Du är efter priset Vadär det? "Han plockade upp lådan och studerade tillbaka." En glöd-in-the-darkbläckfisk! Har du fått ut av det ännu? "Han lutar lådan, vinklasmå färgade bollar av spannmål för att se botten, och nästan spilladem på bordsskivan. "Här är det!" Han släpade ut lite gräddvit,glitter-stänkte bläckfisk, tre inches lång och gjord av gummi plast.
		-- James P. Blaylock, "The Last Coin"

%
Jag fick en antydan om vad som komma när jag hörde min chef klagande, "Theböcker görs och vi fortfarande inte har en författare! Jag måste underteckna någoni dag!på temat läroböcker
		-- Tamim Ansary, "Edutopia Magazine, Issue 2, November 2004"

%
