"Du vet, naturligtvis, att Tasmanians, som aldrig begått äktenskapsbrott, ärnu utdöda. "
		-- M. Somerset Maugham

%
"Om det inte är trasigt, laga det inte."
		-- Bert Lantz

%
"Den charm äktenskapet är att det gör ett liv av bedrägeri en nödvändighet."
		-- Oscar Wilde

%
"Gud är en komiker som spelar för en publik alltför rädda för att skratta."
		-- Voltaire

%
"IBM använder vad jag vill kalla" hole-in-the-marken tekniken "att förstöra konkurrensen ..... IBM gräver ett stort hål imarken och täcker den med löv. Det sätter sedan en stor pottAV GULD i närheten. Då ger samtalet "Hej, titta på alladetta guld, kom hit snabbt. " Så snart konkurrentnärmar potten, faller han i gropen "
		-- John C. Dvorak

%
"Det finns saker som är så allvarliga att du bara kan skämta om dem"
		-- Heisenberg

%
"Det tar alla typer av in och ut-dörr skolgång att få anpassadtill min typ av lurar "
		-- R. Frost

%
"Förbrylla dessa förfäder .... De har stulit våra bästa idéer!"
		-- Ben Jonson

%
Och du skall äta det som korn kakor och du skall baka det med gödsel somgår ut människan, i sin syn ... Sedan han [Herren!] sade till mig, Lo, jaghar gett dig ko dynga för människoträck, och du skall bereda bröddärtill.[Hes. 4: 12-15 (KJV)]
		-- Ben Jonson

%
Jag har skalat bort min klänning; måste jag sätta på den igen? Jag har tvättat mina fötter;måste jag jord dem igen?När min älskade gled handen genom spärren hål, min mage rörsinom mig [mina tarmar flyttades för honom (KJV)].När jag uppstod att öppna för min vän, mina händer dröp av myrra; vätskanmyrra från mina fingrar körde över knoppar av bulten. Med mina egna händer Iöppnas för min kärlek, men min kärlek hade vänt sig bort och gått; mitt hjärta sjönk närHan vände ryggen. Jag sökte honom men jag hittade inte honom, kallade jag honom men hansvarade inte.Väktare, gå rundor i staden, mötte mig; De slog mig och  sårade mig; väktare på väggarna tog bort min mantel.[Visan 5: 3-7 (NEB)]
		-- Ben Jonson

%
Hur vacker är dina fötter med skor, O prins dotter! lederna thylår är som juveler, arbetet i händerna på en slug arbetare. din navelär en rundad skål, som wanteth inte sprit: din buk är som en högvete satte igång med liljor.Din barm är som två unga rosor som är tvillingar.[Visan 7: 1-3 (KJV)]
		-- Ben Jonson

%
Så vackert, hur förtroll du är, min älskade, dotter till läckerheter!Du är ståtlig som en palm, och dina bröst är kluster av datum.Jag sa, "Jag kommer att klättra upp i handflatan att förstå sina ormbunksblad." Kan jag hittabröst som kluster av druvor på vinstockar, doften av din andedräkt somaprikoser och dina viskningar som kryddat vin flyter smidigt att välkomna minsmekningar, glida ner genom läppar och tänder.[Visan 7: 6-9 (NEB)]
		-- Ben Jonson

%
Bär mig som ett sigill på ditt hjärta, som ett sigill vid din arm; Ty kärleken är starksom döden, passion grym som graven; det flammar upp som flammande eld, hårdareän någon flamma.[Visan 8: 6 (NEB)]
		-- Ben Jonson

%
Men Rab-Sake sade till dem, min herre har sänt mig till din herre, ochdig, att tala dessa ord? Har han inte skickade mig till de män som sitter påvägg, så att de kan äta sin egen träck och dricka sitt eget piss med dig?[2 Kings 18:27 (KJV)]
		-- Ben Jonson

%
När HERREN, din gudar har satt dig i det land du ska ockupera, ochdrivas ut många otrogna innan du ... du är att skära ner dem och utrotadem. Du ska inte göra någon kompromiss med dem eller visa dem någon nåd.[Mos. 7: 1 (KJV)]
		-- Ben Jonson

%
Jag tänkte bara på något roligt ... din mamma.
		-- Cheech Marin

%
I början var jag gjort. Jag frågade inte göras. Ingen har hörtmed mig eller anses mina känslor i denna fråga. Men om det tog någradagslända till vissa blyg människor som de på måfå pranced väggenom livets sorgliga djungel, då blir det så.- Marvin Paranoid Android, från Douglas Adams Hitchiker Rens guide tillGalaxy Radio Skript
		-- Cheech Marin

%
Du kommer att lyckas i ditt arbete.
		-- Cheech Marin

%
Livslängden för en repa man är alltid intensiv.
		-- Cheech Marin

%
Om du inte är försiktig, kommer du att fånga något.
		-- Cheech Marin

%
Det är det om personer som tror att de hatar datorer. Vad deverkligen hatar är usel programmerare.
		-- Larry Niven and Jerry Pournelle in "Oath of Fealty"

%
Vart du än går ... Det är du.
		-- Buckaroo Banzai

%
Livet i naturtillståndet är ensam, dålig, otäckt, djuriskt, och kort.
		-- Thomas Hobbes, Leviathan

%
Oskicklighet dikterar ekonomin i stil.
		-- Joey Ramone

%
Ingen är lämplig att lita med kraft. ... Ingen. ... Varje människa som har levtalls känner till dårskaper och ondska han är kapabel till. ... Och om han görvet det, vet han också att varken han eller någon borde fåbesluta en enda människa öde.
		-- C. P. Snow, The Light and the Dark

%
Framgångsrik och lycklig brott kallas förtjänst.
		-- Seneca

%
När vi hoppade in Sicilien, blev enheterna separeras, och jag kunde inte hittanågon. Så småningom jag snubblat över två överstar, en stor, tre kaptener,två löjtnanter och en rifleman, och vi säkrade bron. Aldrig ihistoria av krig har så få letts av så många.
		-- General James Gavin

%
Det enda som krävs för en triumf för det onda är att goda män att göra ingenting.
		-- Edmund Burke

%
Du kan ringa mig av mitt namn, Wirth, eller min värde, Worth.
		-- Nicklaus Wirth

%
Ge en man en fisk, och du matar honom för en dag.Lär en man att fiska, och han kommer att bjuda in sig själv på middag.
		-- Calvin Keegan

%
Förutsägelse är mycket svårt, särskilt när det gäller framtiden.
		-- Niels Bohr

%
Datorn kan inte berätta den känslomässiga historia. Det kan ge dig den exaktamatematisk design, men vad som saknas är ögonbrynen.
		-- Frank Zappa

%
Saker och ting är inte så enkla som de verkar vid första.
		-- Edward Thorp

%
Huvudsaken är att spela själv. Jag svär att girighet för pengarna har ingentingatt göra med det, även om himlen vet jag verkligen i behov av pengar.
		-- Feodor Dostoyevsky

%
Det är säkerligen en stor olycka för en människa att ha några tvångstankar.
		-- Robert Bly

%
Maskiner tar mig på sängen med stor frekvens.
		-- Alan Turing

%
Osäker förmögenhet noggrant behärskas av det egna kapitalet i beräkningen.
		-- Blaise Pascal

%
Efter Goliats nederlag, jättar upphörde att befalla respekt.
		-- Freeman Dyson

%
Det finns två sätt att konstruera en programvara design. Ett sätt är att göradet så enkelt att det inte är självfallet inga brister och den andra är attgöra det så komplicerat att det inte finns några uppenbara brister.
		-- Charles Anthony Richard Hoare

%
Låt inte detta språk (Ada) i sitt nuvarande tillstånd för att användas iapplikationer där tillförlitlighet är kritiska, dvs kärnkraftverk,kryssningsmissiler, system för tidig varning, anti-ballistiska missilförsvarsystem. Nästa raket för att gå vilse som ett resultat av ett programmeringsspråkfel kan inte vara ett förberedande rymdraket på en ofarlig resa till Venus:Det kan vara en kärnstridsspetsar exploderar över en av våra städer. en opålitligprogrammeringsspråk genere opålitliga program utgör en mycketstörre risk för vår miljö och vårt samhälle än osäkra bilar, giftigbekämpningsmedel, eller olyckor vid kärnkraftverk.
		-- C. A. R. Hoare

%
Utan kaffe han inte kunde arbeta, eller åtminstone han inte kunde har arbetat isätt han gjorde. Förutom papper och pennor, tog han med sig överallt som enoumbärlig artikel av utrustning kaffemaskinen, som var mindreviktigare för honom än hans bord eller sin vita dräkt.
		-- Stefan Zweigs, Biography of Balzac

%
"Det var havsrätts, sa de. Civilization slutar vid vattenlinjen.Utöver detta, vi alla in i livsmedelskedjan, och inte alltid rätt på toppen. "
		-- Hunter S. Thompson

%
I ynklig, sidiga, förbindelse boxed form som flödesschemat haridag utarbetats, det har visat sig vara värdelös som ett designverktyg -programmerare rita flödesscheman efter, inte före, skriver de program debeskriva.
		-- Fred Brooks, Jr.

%
Den så kallade "stationära metafor" av dagens arbetsstationer är istället en"Flygplan-sits" metafor. Den som har blandas en mantel full av papper medansitter mellan två portly passagerare kommer att känna igen skillnaden - en kanse bara en mycket få saker på en gång.
		-- Fred Brooks, Jr.

%
... När anfall av kreativitet köra stark, mer än en programmerare eller författare harvarit kända för att överge skrivbordet för rymligare golvet.
		-- Fred Brooks, Jr.

%
En liten tillbakablickande visar att även om många fina, användbara mjukvarusystemhar utformats av utskotten och byggdes som en del av flera delar projekt,dessa mjukvarusystem som har glada passionerade fans är de som ärprodukter från en eller ett fåtal utforma sinnen, stora designers. Överväga Unix,APL, Pascal, Modula, Smalltalk-gränssnittet, även Fortran; och kontras demmed Cobol, PL / I, Algol, MVS / 370, och MS-DOS.
		-- Fred Brooks, Jr.

%
... Hårdvara framsteg är så snabb. Ingen annan teknik sedancivilisation började har sett sex storleksordningar i prestations prisvinna på 30 år.
		-- Fred Brooks, Jr.

%
Programenheter är mer komplexa för sin storlek än kanske någon annan människakonstruera eftersom det inte finns två delar som är likadana. Om de är, gör vi tvåliknande delar i en subrutin - öppen eller stängd. I detta avseende, mjukvarasystem skiljer sig i grunden från datorer, byggnader eller bilar, därupprepade element i överflöd.
		-- Fred Brooks, Jr.

%
Digitala datorer är själva mer komplex än de flesta saker folk bygga:De har ett mycket stort antal stater. Detta gör att utforma, beskriver,och testa dem hårt. Mjukvarusystem har order-of-magnitud flera staterän datorer gör.
		-- Fred Brooks, Jr.

%
Komplexiteten av programvara är en viktig egenskap, inte ett misstag en.Därför, beskrivningar av en programvara enhet som abstrakt bort dess komplexitetofta abstrakt bort dess väsen.
		-- Fred Brooks, Jr.

%
Einstein menade att det måste förenklas förklaringar av naturen, eftersomGud är inte nyckfull eller godtycklig. Ingen sådan tro tröstar programvaraningenjör.
		-- Fred Brooks, Jr.

%
Med undantag för 75% av kvinnorna, alla i hela världen vill ha sex.
		-- Ellyn Mustard

%
Sambandet mellan det språk som tror att vi / program och de problemoch lösningar som vi kan föreställa oss är mycket nära. Av denna anledning begränsandespråkfunktioner med avsikten att eliminera programmerare fel är i bästa fallfarlig.
		-- Bjarne Stroustrup in "The C++ Programming Language"

%
Det enda sättet att lära sig ett nytt programmeringsspråk är genom att skriva program i den.
		-- Brian Kernighan

%
Perfektion uppnås endast på väg att kollapsa.
		-- C. N. Parkinson

%
Där går man,Hålla så cool som du kan.Det riles dem att tro att du uppfattar webben de väver.Fortsätter att vara gratis!
		-- C. N. Parkinson

%
Bingo, bensinstation, hamburgare med en sida för flygbuller,och du kommer att Gary, Indiana. - Jessie i filmen "Greaser palats"
		-- C. N. Parkinson

%
I hopp om att godhet är inte teologiskt ljud. - Jordnötter nötter~~POS=HEADCOMP
		-- C. N. Parkinson

%
Polisen upp dina oönskade rundor och frags. Låt inte ingenting för dinks.
		-- Willem Dafoe in "Platoon"

%
"Hela mitt liv har jag velat vara någon, jag antar att jag borde ha varit mer specifik."
		-- Jane Wagner

%
"Alla medel tillräckligt kraftfull för att förlänga människans räckvidd är tillräckligt kraftfull för att störtahans värld. För att få mediets magi för att arbeta för sina mål snarare änmot dem är att uppnå och skrivkunnighet. "
		-- Alan Kay, "Computer Software", Scientific American, September 1984

%
"Datakunskap är en kontakt med aktiviteten att beräkna tillräckligt djup för attgöra beräknings motsvarande läsa och skriva flytande och trevlig.Som i alla konst, måste en romans med materialet är på god väg. OmVi värdesätter livslångt lärande av konst och bokstäver som en språngbräda förpersonlig och samhällelig utveckling, bör alla mindre ansträngning spenderas för att göra datoren del av våra liv? "
		-- Alan Kay, "Computer Software", Scientific American, September 1984

%
"De största krigare är de som kämpar för fred."
		-- Holly Near

%
"Oavsett var du går, där är du ..."
		-- Buckaroo Banzai

%
Inkräktare kommer att skjutas. Överlevande kommer att åtalas.
		-- Buckaroo Banzai

%
Inkräktare kommer att skjutas. Överlevande kommer att skjutas IGEN!
		-- Buckaroo Banzai

%
"Jag växer äldre, men inte upp."
		-- Jimmy Buffett

%
Forskarna kommer att studera din hjärna att lära mer om din avlägsen kusin, man.
		-- Jimmy Buffett

%
"Jag hatar klåda. Men jag har inget emot svullnad."- Nya buzz fras som "Var är nötköttet?" att David Letterman försöker   att få alla att börja säga
		-- Jimmy Buffett

%
Din egen lycka kan variera.
		-- Jimmy Buffett

%
"Oh dear, jag tror att du hittar verklighetens på blinkar igen."
		-- Marvin The Paranoid Android

%
"Skicka advokater, vapen och pengar ..."
		-- Lyrics from a Warren Zevon song

%
"Jag går på att arbeta för samma anledning en höna fortsätter lägger ägg."
		-- H. L. Mencken

%
"Kom ihåg att information är inte kunskap, Kunskap är inte visdom;Visdom är inte sanning; Sanningen är inte skönhet, Skönhet är inte kärlek;Kärlek är inte musik; Musik är den bästa. "- Frank Zappa
		-- H. L. Mencken

%
Jag kan inte köra 55.
		-- H. L. Mencken

%
"Och de berättade vad de ville ... Var ett ljud som skulle kunna döda någon-en, från ett avstånd. "- Kate Bush
		-- H. L. Mencken

%
"Mot bakgrund av entropi och intet, du slags måste låtsas att det är intedär om du vill fortsätta skriva bra kod. "- Karl Lehenbauer
		-- H. L. Mencken

%
Märken? Vi behöver inte några stinkande märken.
		-- H. L. Mencken

%
Jag kan inte köra 55.Jag ser fram emot att inte kunna köra 65, heller.
		-- H. L. Mencken

%
Tack och lov en miljon miljarder gånger du bor i Texas.
		-- H. L. Mencken

%
"Kan du programmera?" "Ja, jag är skrivkunnig, om det är vad du menar!"
		-- H. L. Mencken

%
Inga användar servicable delar inuti. Se till kvalificerad servicepersonal.
		-- H. L. Mencken

%
I hjärtat av vetenskap är en viktig spänning mellan två till synesmotsägelsefulla attityder - en öppenhet för nya idéer, oavsett hur bisarraeller bakvända de kan vara, och mest hänsynslösa skeptiska granskningav alla idéer, gamla och nya. Detta är hur djupt sanningar sållas från djupdumheter. Naturligtvis, forskare göra misstag för att försöka förståvärlden, men det finns en inbyggd felkorrigerande mekanism: Den kollektivaföretag i kreativt tänkande och skeptiska tänkande tillsammans hållerfält på rätt spår.
		-- Carl Sagan, "The Fine Art of Baloney Detection," Parade, February 1, 1987

%
En av de sorgligaste lärdom av historien är här: Om vi ​​har bamboozledtillräckligt länge, tenderar vi att avvisa alla bevis på Bamboozle. Vi är intelängre är intresserad av att ta reda på sanningen. Den Bamboozle har fångatoss. det är helt enkelt alltför smärtsamt att erkänna - även för oss själva - attVi har varit så godtrogna. (Så gamla Bamboozles tenderar att kvarstå somnya Bamboozles stiga.)
		-- Carl Sagan, "The Fine Art of Baloney Detection," Parade, February 1, 1987

%
Beträffande astral projektion, Woody Allen skrev en gång, "Detta är inte ett dåligt sättatt resa, även om det är oftast en halvtimme vänta för bagage. "
		-- Carl Sagan, "The Fine Art of Baloney Detection," Parade, February 1, 1987

%
Oförmågan att dra nytta av återkoppling verkar vara den primära orsaken tillpseudovetenskap. Pseudo behålla sin tro och ignorera eller förvrängamotsägelsefulla bevis snarare än ändra eller avvisa en bristfällig teori. Därför attav deras starka fördomar, de verkar sakna självkorrigerande mekanismerforskare måste använda i sitt arbete.
		-- Thomas L. Creed, "The Skeptical Inquirer," Summer 1987

%
Att hitta enstaka halm sanning översköljs i en stor ocean av förvirring ochBamboozle kräver intelligens, vaksamhet, engagemang och mod. Men om viinte utövar dessa tuffa tankevanor, kan vi inte hoppas på att lösa de verkligtallvarliga problem som möter oss - och vi riskerar att bli en nation av rotskott, uppslåss av nästa charlatan som kommer tillsammans.
		-- Carl Sagan, "The Fine Art of Baloney Detection," Parade, February 1, 1987

%
Inte underskatta värdet av tryckta rapporterna för felsökning.
		-- Carl Sagan, "The Fine Art of Baloney Detection," Parade, February 1, 1987

%
Inte underskatta värdet av tryckta rapporterna för felsökning.Har inte estetiska kramper när du använder dem, heller.
		-- Carl Sagan, "The Fine Art of Baloney Detection," Parade, February 1, 1987

%
Eftersom systemet kommer upp, kommer komponentbyggare från tid till annan visasbärande heta nya versioner av sina pjäser - snabbare, mindre, mer kompletta,eller förmodat mindre buggy. Ersättandet av en arbetande komponent med en nyversionen kräver samma systematiska testförfarande som lägger till en nykomponent gör, även om det skulle kräva mindre tid för mer komplett ocheffektiva testfall vanligtvis tillgängliga.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Varje teambuilding annan komponent har använt den senaste testadeversion av det integrerade systemet som en provbänk för felsökning sin pjäs. DerasArbetet kommer att ställa tillbaka genom att ha att provbänk förändring under dem. Naturligtvis är detmåste. Men förändringarna måste vara kvantiserade. Då varje användare har perioder avproduktiv stabilitet, avbruten av skurar av testbädd förändring. detta verkaratt vara mycket mindre störande än en konstant porlande och darrande.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Begrepps integritet i sin tur kräver att konstruktionen måste utgå från ensinne, eller från ett mycket litet antal enas resonans sinnen.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Det är en mycket ödmjuka upplevelse att göra en mångmiljondollar misstag, men detär också mycket minnesvärd. Jag minns tydligt natten vi beslutat hur man organiserarsjälva skrivandet av externa specifikationer för OS / 360. Chef förarkitektur, chef för genomförandet styrprogram, och jag vartröska ut planen, schema och ansvarsfördelning.Arkitekturen chef hade 10 goda män. Han hävdade att de kunde skrivaspecifikationer och gör det rätt. Det skulle ta tio månader, tre merän schemat tillåtet.Kontrollprogrammet chef hade 150 män. Han hävdade att de kunde förberedaspecifikationerna, med arkitekturen laget samordnande; det skulle varavälgjord och praktisk, och han kunde göra det på schemat. Dessutom, omarkitekturen laget gjorde det, skulle hans 150 män sitta tråkigt sina tummari tio månader.Till detta svarade arkitektur chefen att om jag gav styrprogrammetlaget ansvar, skulle resultatet i själva verket inte vara på gång, men skulleockså vara tre månader för sent, och mycket lägre kvalitet. Jag gjorde, och det var. hanvar rätt på båda dessa punkter. Dessutom bristen på begrepps integritet gjortsystemet betydligt mer kostsamt att bygga och förändring, och jag skulle uppskatta att detlagt ett år till felsökning tid.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Anledningen ESP, till exempel, anses inte vara en livskraftig ämne i dagenspsykologi är helt enkelt att utredningen inte har visat sig vara fruktbart ... Eftermer än 70 års studier, det fortfarande inte finns ett exempel på en ESPfenomen som är repliker under kontrollerade förhållanden. Denna enkla mengrundläggande vetenskapliga kriteriet inte har uppfyllts trots dussintals studierunder många decennier ... Det är av detta skäl att ämnet är nu litenintresse för psykologi ... Kort sagt, det finns ingen visat fenomen sombehöver förklaring.
		-- Keith E. Stanovich, "How to Think Straight About Psychology", pp. 160-161

%
Utvecklingen av den mänskliga rasen kommer inte ske i tiotusenår av tama djur, men i miljoner år av vilda djur, eftersom manär och kommer alltid att vara ett vilt djur.
		-- Charles Galton Darwin

%
Naturligt urval kommer ingen roll snart, inte någonstans så mycket som medvetet val.Vi kommer att civilisera och förändra oss för att passa våra idéer om vad vi kan vara.Inom en mer mänsklig livslängd, kommer vi att ha ändrat oss oigenkännlighet.
		-- Greg Bear

%
"Jesus kan älska dig, men jag tror att du är skräp insvept i huden."
		-- Michael O'Donohugh

%
... Men hans uppfinning fungerade utmärkt - hans teori var en kruka av avloppsvatten frånbörjan till slut. - Vernor Vinge, "The Peace War"
		-- Michael O'Donohugh

%
"Det är som deja vu igen." - Yogi Berra
		-- Michael O'Donohugh

%
Det sista man vet att konstruera ett verk är vad man ska sätta först.
		-- Blaise Pascal

%
"Var ska jag börja, vänligen Ers Majestät?" han frågade. "Börja från början"kungen sade, allvarligt, "och gå på tills du kommer till slutet. sedan stoppa"Alice i Underlandet, Lewis Carroll
		-- Blaise Pascal

%
En bit av äkta historia är en sak så sällsynt som att alltid vara värdefull.
		-- Thomas Jefferson

%
Att vara vaken är att vara vid liv. - Henry David Thoreau, i "Walden"
		-- Thomas Jefferson

%
En person med en klocka vet vilken tid det är; en person med två klockor äraldrig säker. Ordspråk
		-- Thomas Jefferson

%
Du ser men inte observera.Sir Arthur Conan Doyle, i "The Memoirs of Sherlock Holmes"
		-- Thomas Jefferson

%
Ett gräl snabbt avvecklas när övergiven av en part; det finns ingen kampsåvida det finnas två. - Seneca
		-- Thomas Jefferson

%
Ingenting någonsin blir verklighet tills det upplevs - även ett ordspråk är ingen ordspråktill dig tills ditt liv har illustrerat det. - John Keats
		-- Thomas Jefferson

%
Fancy är verkligen inget annat än en form av minne frigjord från beställningenav tid och rum. - Samuel Taylor Coleridge
		-- Thomas Jefferson

%
Vad vi förväntar oss sällan inträffar; vad vi minst anar i allmänhet händer.
		-- Bengamin Disraeli

%
Ingenting i progression kan vila på sin ursprungliga plan. Vi kan lika gärna tänka pågunga en vuxen man i vaggan för ett spädbarn. - Edmund Burke
		-- Bengamin Disraeli

%
För varje problem finns det en lösning som är enkel, snygg, och fel.
		-- H. L. Mencken

%
Säg inte hur hårt du arbetar. Säg mig hur mycket du får gjort.
		-- James J. Ling

%
En vän i livet är mycket; två är många; tre är knappast möjligt.Vänskap behöver en viss parallellitet i livet, en gemenskap av tanken,en rivalitet av mål. - Henry Brook Adams
		-- James J. Ling

%
Kom ihåg digAy, du dålig spöke medan minnet har en sitsI detta distraherad jordklotet. Kom ihåg dig!Ja, från bordet av mitt minneJag ska torka bort alla triviala förtjust poster,Alla sågar av böcker, alla former, alla tryck förbi,Att ungdomar och observation kopieras dit.Hamlet, I: v: 95 William Shakespeare
		-- James J. Ling

%
Självklart kan man dom inte vara bättre än den information som hangrundar det. Ge honom sanningen och han kan fortfarande gå fel när han harchansen att vara rätt, men ger honom inga nyheter eller presentera honom endast med förvrängdoch ofullständiga uppgifter, med okunniga, slarvig eller partisk rapportering, med propagandaoch avsiktliga lögner och du förstöra hans hela resonemang processer, ochgöra honom något mindre än en människa.
		-- Arthur Hays Sulzberger

%
Varje ärlig samtal, varje promenad i livet, har sin egen elit, sin egen aristokratibaserad på spetskompetens prestanda. - James Bryant Conant
		-- Arthur Hays Sulzberger

%
Du kan observera en hel del bara genom att titta på. - Yogi Berra
		-- Arthur Hays Sulzberger

%
Om närvaron av elektricitet kan synliggöras i någon del av en krets, jagser ingen anledning till varför intelligens inte kan överföras omedelbart efterelektricitet. - Samuel F. B. Morse
		-- Arthur Hays Sulzberger

%
"Mr Watson, kom hit, jag vill ha dig." - Alexander Graham Bell
		-- Arthur Hays Sulzberger

%
Det är för närvarande ett problem att få tillgång till gigabit via punybaud.
		-- J. C. R. Licklider

%
Det är viktigt att notera att troligen ingen stor operativsystem med dagenskonstruktionsteknik kan motstå en bestämd och väl samordnat angrepp,och att de flesta sådana dokumenterade genomföringar har varit förvånansvärt lätt.- B. Hebbard "A Penetration Analys av Michigan terminalsystem",Operativsystem Review, Vol. 14, nr 1, juni 1980, sid. 7-20
		-- J. C. R. Licklider

%
En rätt är inte vad någon ger dig; det är vad ingen kan ta ifrån dig.
		-- Ramsey Clark

%
Priset man betalar för att uppnå något yrke, eller ringa, är en intimkunskap om sitt fula sida. - James Baldwin
		-- Ramsey Clark

%
Litet är vackert.
		-- Ramsey Clark

%
... Den ökade produktiviteten främjas av en vänlig miljö och kvalitetverktyg är avgörande för att möta de ständigt ökande kraven på programvara.
		-- M. D. McIlroy, E. N. Pinson and B. A. Tague

%
Det är inte bäst att byta hästar när de korsar floden.
		-- Abraham Lincoln

%
Speglar bör återspegla lite innan man kastar upp bilder.
		-- Jean Cocteau

%
Antag för ett ögonblick att bilindustrin hade utvecklats på sammatakt som datorer och under samma period: hur mycket billigare och effektivareskulle de nuvarande modellerna vara? Om du inte redan har hört analogtSvaret är splittring. Idag skulle du kunna köpa en Rolls-Royce för $ 2,75,det skulle göra tre miljoner miles till gallon, och det skulle ge tillräckligtkraft för att driva Queen Elizabeth II. Och om du var intresserade avminiatyrisering, kan du placera ett halvt dussin av dem på ett knappnålshuvud.
		-- Christopher Evans

%
I framtiden kommer du att få datorer som priser i frukostflingor.Du kastar ut dem eftersom ditt hus kommer att kantas dem.
		-- Robert Lucky

%
Få tag i bärbara egendom. - Charles Dickens, "Stora förväntningar"
		-- Robert Lucky

%
Sammantaget är filosofin att angripa tillgänglighet problemet från tvåkompletterande riktningar: att minska antalet mjukvaru fel genomrigorösa tester för att driva system, och för att minska effekten avåterstående fel genom att för återvinning av dem. En intressant fotnottill denna konstruktion är att nu kan vanligtvis betraktas som ett systemfel att vararesultatet av två program fel: den första, i det program som startadeproblem; den andra, i återhämtningen rutin som inte kunde skyddasystem. - A. L. Scherr, "Functional struktur IBM Virtual Storage RörelseSystem, del II: OS / VS-2 Begrepp och filosofier, "IBM Systems Journal,Vol. 12, nr 4, 1973, sid. 382-400
		-- Robert Lucky

%
Hur många hårdvara killar tar det att byta en glödlampa?"Jo diagnostiken säger att det är bra kompis, så det är ett programvaruproblem."
		-- Charles Babbage, Passage from the Life of a Philosopher

%
"Försök inte outweird mig, tre ögon. Jag får konstigare saker än du gratismed min frukostflingor. "
		-- Zaphod Beeblebrox in "Hitchiker's Guide to the Galaxy"

%
Okompenserad övertid? Säg bara nej.
		-- Zaphod Beeblebrox in "Hitchiker's Guide to the Galaxy"

%
Koffeinfritt kaffe? Säg bara nej.
		-- Zaphod Beeblebrox in "Hitchiker's Guide to the Galaxy"

%
"Showbusiness är precis som high school, förutom att du får betalt."
		-- Martin Mull

%
"Detta är inte en hjärnoperation, det är bara tv."
		-- David Letterman

%
"Moral är en sak. Betyg är allt."
		-- A Network 23 executive on "Max Headroom"

%
Lev fritt eller dö.
		-- A Network 23 executive on "Max Headroom"

%
"... Om kyrkan sätta på halva tiden på girighet som det gör på lust, detta skulle vara en bättre värld. "- Garrison Keillor," Lake Wobegon Days "
		-- A Network 23 executive on "Max Headroom"

%
Utanför en hund, en bok man bästa vän. Inuti en hund, är det ocksåmörk att läsa.
		-- A Network 23 executive on "Max Headroom"

%
"Förmodligen det bästa operativsystemet i världen är [operativsystem] gjorts för PDP-11 av Bell Laboratories. "- Ted Nelson, oktober 1977
		-- A Network 23 executive on "Max Headroom"

%
"Alla dessa svarta människor skruva upp min demokrati." - Ian Smith
		-- A Network 23 executive on "Max Headroom"

%
Använd Force, Luke.
		-- A Network 23 executive on "Max Headroom"

%
Jag har en dålig känsla om detta.
		-- A Network 23 executive on "Max Headroom"

%
Befogenhet att förstöra en planet är obetydlig i jämförelse med kraften ikraften.
		-- Darth Vader

%
När jag lämnade dig, var jag men eleven. Nu är jag befälhavaren.
		-- Darth Vader

%
"Ja, ja, ja! Tja om det är inte fett stinkande bocken Billy Boy iförgifta! Hur du, du globby flaska billig stinkande chip olja? Kommaoch få en i yarbles, om ya har någon yarble, ya eunuck gelé du! "
		-- Alex in "Clockwork Orange"

%
"Det fanns inget jag hatade mer än att se en smutsig gammal Drunkie, ett tjutandebort på söner sin far och går blurp Blurp mellan som om det voreen snuskig gammal orkester i sin stinkande ruttna tarmar. Jag kunde aldrig stå tillse någon sådär, särskilt när de var gamla som denna var. "
		-- Alex in "Clockwork Orange"

%
186.000 Miles per sekund. Det är inte bara en bra idé. Det är lagen.
		-- Alex in "Clockwork Orange"

%
Dumhet, som dygd, är sin egen belöning.
		-- Alex in "Clockwork Orange"

%
Gee, Toto, jag tror inte att vi är i Kansas anymore.
		-- Alex in "Clockwork Orange"

%
Barn börjar genom att älska sina föräldrar. Efter en tid som de bedömer dem. Sällan,om någonsin, de förlåter dem.
		-- Oscar Wilde

%
Enda tasking: Just Say Nej
		-- Oscar Wilde

%
"Fånga en våg och du sitter på toppen av världen."
		-- The Beach Boys

%
"Bond återspeglas att goda amerikaner var fina människor och att de flesta av demtycktes komma från Texas. "
		-- Ian Fleming, "Casino Royale"

%
"Jag tror att skräp är den viktigaste manifestation av kultur vi har i minlivstid."
		-- Johnny Legend

%
Med en räkning finns några 700 forskare med respektabla akademiska meriter(Av totalt 480.000 amerikanska jord och livs forskare) som ger trovärdighetskapandet-vetenskap, den allmänna teorin att komplexa livsformer inte utvecklasmen verkade "abrupt".
		-- Newsweek, June 29, 1987, pg. 23

%
Även om du kan lura folk om en produkt genom vilseledande uppgifter,förr eller senare kommer produkten att tala för sig själv.
		-- Hajime Karatsu

%
För att lyckas i något företag, måste man vara långlivade och patient.Även om man måste köra vissa risker, måste man vara modig och stark nog attmöta och övervinna besvärliga utmaningar för att upprätthålla ett framgångsrikt företag ipå lång sikt. Jag kan inte låta bli att säga att amerikaner saknar detta nödvändigtutmanande anda idag.
		-- Hajime Karatsu

%
Minnen av du påminner mig om dig.
		-- Karl Lehenbauer

%
Liv. Prata inte med mig om livet.
		-- Marvin the Paranoid Android

%
En klar skiva kan du söka evigt.
		-- Marvin the Paranoid Android

%
Världen går mot sitt slut - spara buffertar!
		-- Marvin the Paranoid Android

%
grep mig inga mönster och jag ska säga dig inga linjer.
		-- Marvin the Paranoid Android

%
Det är ditt öde.
		-- Darth Vader

%
Lucas religioner och antika vapen är ingen ersättning för en bra blaster pådin sida.
		-- Han Solo

%
Hur många QA ingenjörer tar det att skruva i en glödlampa?3: 1 för att skruva in den och två att säga "jag sa" när det inte fungerar.
		-- Han Solo

%
Hur många NASA chefer tar det att skruva i en glödlampa?"Det är ett känt problem ... inte oroa sig för det."
		-- Han Solo

%
Att vara är att programmera.
		-- Han Solo

%
Till programmet är att vara.
		-- Han Solo

%
Jag programmerar, därför är jag.
		-- Han Solo

%
Människor är mycket flexibla och lära sig att anpassa sig till främmandeomgivning - de kan bli vana vid att läsa Lisp ochFortran program, till exempel.
		-- Leon Sterling and Ehud Shapiro, Art of Prolog, MIT Press

%
"Jag är din densitet."
		-- George McFly in "Back to the Future"

%
"Så varför inte du göra som ett träd, och få outta här."
		-- Biff in "Back to the Future"

%
"Falling in love gör rökning potten hela dagen ser ut som den ultimata återhållsamhet."
		-- Dave Sim, author of Cerebrus.

%
Guds existens innebär en kränkning av orsakssamband.
		-- Dave Sim, author of Cerebrus.

%
"Jag kan kid runt om droger, men egentligen, jag tar dem på allvar."
		-- Doctor Graper

%
Operativsystemet programvara är program som dirigerar alla grundläggandefunktionerna hos en dator.
		-- The Wall Street Journal, Tuesday, September 15, 1987, page 40

%
Jag svär trohet till flaggani Amerikas förenta stateroch till republiken som den står för,en nation,odelbar,med frihetoch rättvisa för alla.
		-- Francis Bellamy, 1892

%
Folk tror att min vän George är konstigt eftersom han bär polisonger ... bakom hansöron. Jag tror att han är konstigt eftersom han bär löständer ... med hängslen på dem.
		-- Steven Wright

%
Min bror skickade mig ett vykort häromdagen med denna stora satellitbildhela jorden på den. På baksidan det sade: "Önskar du var här".
		-- Steven Wright

%
Du kan inte få allt ... var skulle du placera den?
		-- Steven Wright

%
Jag spelade poker häromkvällen ... med tarotkort. Jag fick en kåk och4 personer dog.
		-- Steven Wright

%
Du vet den där känslan när du lutade sig tillbaka på en pall och det börjar att tippaöver? Tja, det är hur jag känner hela tiden.
		-- Steven Wright

%
Jag kom hem den andra natten och försökte öppna dörren med mina bilnycklar ... ochbyggnaden startas. Så jag tog ut för en enhet. En polis drog mig överför fortkörning. Han frågade mig där jag bor ... "Här".
		-- Steven Wright

%
"Leva eller dö, jag ska göra en miljon."
		-- Reebus Kneebus, before his jump to the center of the earth, Firesign Theater

%
Den typiska sidlayout program är inget annat än en elektroniskljusbord för skärning och klistra dokument.
		-- Reebus Kneebus, before his jump to the center of the earth, Firesign Theater

%
Det finns buggar och sedan finns det buggar. Och sedan finns det buggar.
		-- Karl Lehenbauer

%
Min dator kan slå upp datorn.
		-- Karl Lehenbauer

%
Döda Ugly processorarkitekturer
		-- Karl Lehenbauer

%
Döda Ful Radio
		-- Frank Zappa

%
"Säg bara nej." - Nancy Reagan"Nej." - Ronald Reagan
		-- Frank Zappa

%
Jag tror att en del av det som driver vetenskapen är törst efter att undra. Det är enmycket kraftfulla känslor. Alla barn känner det. I en första klass klassrumalla känner det; i en tolfte klass klassrum nästan ingen känner det, elleråtminstone erkänner det. Något händer mellan första och tolfte klass,och det är inte bara puberteten. Inte bara de skolor och media inte undervisamycket skepsis, det finns också lite uppmuntran av denna omrörda känslaav förundran. Vetenskap och pseudovetenskap både väcka den känslan. Fattigpopulariseringar vetenskapens inrätta en ekologisk nisch för pseudovetenskap.
		-- Carl Sagan, The Burden Of Skepticism, The Skeptical Inquirer, Vol. 12, Fall 87

%
Om vetenskapen förklarades för en vanlig människa på ett sätt som är tillgängligtoch spännande, skulle det inte finnas något utrymme för pseudovetenskap. Men det finns en sortsav Gresham lag genom vilken i populärkulturen dålig vetenskap driver utbra. Och för detta jag tror att vi måste skylla, första, det vetenskapliga samfundetoss för att inte göra ett bättre jobb popularisera vetenskap, och för det andramedier, som är i detta avseende nästan jämnt fruktansvärda. varje tidningi Amerika har en daglig astrologi kolonn. Hur många har även en gång i veckanastronomi kolonn? Och jag tror att det är också fel utbildningssystem. Vi lär inte ut hur man tänker. Detta är en mycket allvarlig brist somkan även, i en värld riggad med 60.000 kärnvapen, äventyra människorsframtida.
		-- Carl Sagan, The Burden Of Skepticism, The Skeptical Inquirer, Vol. 12, Fall 87

%
"Jag hävdar att det är mycket mer konstigt i vetenskap än i pseudovetenskap. OchFörutom att det mått denna term har någon mening, har vetenskapenytterligare stöd, och det är inte en obetydlig en, för att vara sant.
		-- Carl Sagan, The Burden Of Skepticism, The Skeptical Inquirer, Vol. 12, Fall 87

%
Jag får ofta frågan frågan, "Tror du att det finns utomjordiska intelli-? Gens "Jag ger standard argument - det finns en hel del platser där ute,och använda ordet * miljarder *, och så vidare. Och då säger jag att det skulle vara förvånandetill mig om det inte fanns utomjordisk intelligens, men naturligtvis finns det sommen inga övertygande bevis för det. Och då jag frågade, "Ja, men vad gör duverkligen tror? "Jag säger:" Jag sa ju vad jag tycker egentligen. "" Ja, menVad är din magkänsla? "Men jag försöker att inte tänka med min gut. Egentligen är detokej att reservera dom tills bevisen är i.
		-- Carl Sagan, The Burden Of Skepticism, The Skeptical Inquirer, Vol. 12, Fall 87

%
Stöta bort dem. Stöta bort dem. Förmå dem att avstå från sfäroid.
		-- Indiana University fans' chant for their perennially bad football team

%
Om det fungerar, diagnostiken säger att det är bra.Om det inte fungerar, diagnostiken säger att det är bra.
		-- A proposed addition to rules for realtime programming

%
   Det är antingen genom påverkan av narkotiska potions, varav allaprimitiva folk och raser tala i psalmer, eller genom kraftfull metodav våren, genomträngande med glädje hela naturen, att de dionysiska rörelsernauppstå, vilket i sin intensifiering leda individen att glömma sig självfullständigt. . . .Inte Bara gör bandet mellan människa och människa kommit att smiddaåterigen av den magiska dionysiska rit, men alienerade, fientlig, ellerunderkuvade naturen firar igen hennes försoning med sin förlorade sonen,man.
		-- Fred Nietzsche, The Birth of Tragedy

%
Den karakteristiska egenskapen hos hallucinogener, att upphäva gränserna mellandet upplevande själv och den yttre världen i en extatisk, känslomässig upplevelse,gör det möjligt att med deras hjälp, och efter lämplig intern och externpreparatet ... att framkalla en mystisk upplevelse enligt plan, så att säga ...Jag ser den sanna betydelsen av LSD i möjligheten att ge materiellt biståndtill meditation som syftar till den mystiska upplevelsen av en djupare, omfattandeverklighet. En sådan användning överensstämmer helt med det väsentliga och arbetar karaktärLSD som en helig läkemedel.
		-- Dr. Albert Hoffman, the discoverer of LSD

%
Jag delar tron ​​på många av mina samtida att den andliga krisgenomsyrar alla områden i västra industrisamhället kan endast åtgärdasgenom en förändring i vår syn på världen. Vi måste övergå från materialistiska,dualistiska tro att människor och deras miljö är separat, mot enny medvetenhet om en allomfattande verklighet, som omfamnarupplever ego, en verklighet där människor känner att deras enhet med levandenatur och hela skapelsen.
		-- Dr. Albert Hoffman

%
Avsiktlig provokation av mystisk upplevelse, särskilt genom LSD och tillhörandehallucinogener, i motsats till spontana visionära upplevelser, medförfaror som inte får underskattas. Utövare måste ta hänsynhänsyn till de speciella effekterna av dessa ämnen, nämligen deras förmåga tillpåverka vårt medvetande, den innersta kärnan i vår varelse. HistorienLSD hittills visar tydligt de katastrofala följder som kanuppstå när dess djupa effekt missbedömde och ämnet är felför en glädje drog. Särskilda interna och externa preparat förskottkrävs; med dem, kan en LSD experiment bli en meningsfullerfarenhet.
		-- Dr. Albert Hoffman, the discoverer of LSD

%
Jag tror att om folk skulle lära sig att använda LSD vision framkallande förmågaklokare, under lämpliga förhållanden, i medicinsk praxis och i sambandmed meditation, sedan i framtiden problemet barn kan bli ett konstigtbarn.
		-- Dr. Albert Hoffman, the discoverer of LSD

%
I området för vetenskaplig observation, är tur beviljas endast till dem som ärberedd.
		-- Louis Pasteur

%
core fel - buss dumpade
		-- Louis Pasteur

%
Om präglade folieförseglingen undersjal är trasig eller saknas när köpt, inteanvändning.
		-- Louis Pasteur

%
"Kom hit, baby, jag vill göra en sak med dig."
		-- A Cop, arresting a non-groovy person after the revolution, Firesign Theater

%
"Ahead varp faktor 1"
		-- Captain Kirk

%
   Eldig energi lanced ut, men balkarna slog en immateriell vägg mellanden Gubru och snabbt vända jorden skepp.   "Vatten!" det skrek som läser den spektrala rapport. "En barriär av vattenånga! Ett civiliserat ras kunde inte ha hittat en trick i biblioteket!Ett civiliserat ras kunde inte ha böjde så låg! Ett civiliserat ras skulle inteha..."   Det skrek som Gubru fartyget slog ett moln av drivande snöflingor.
		-- Startide Rising, by David Brin

%
Harrison postulatet:För varje handling finns en likvärdig och motsatt kritik.
		-- Startide Rising, by David Brin

%
Mr Coles Axiom:Summan av intelligens på planeten är en konstant;befolkningen växer.
		-- Startide Rising, by David Brin

%
Felson lag:Att stjäla idéer från en person är plagiat; att stjäla frånmånga är forskning.
		-- Startide Rising, by David Brin

%
... En annan författare igen överens med alla mina generaliseringar, men sade att som eninbiten skeptiker Jag har stängt min sinne för sanningen. Framför allt har jagignorerat bevis för en jord som är sex tusen år gammal. Tja, jaghar inte ignorerat det; Jag ansåg den påstådda bevis och * sedan * förkastade det.Det finns en skillnad, och det är en skillnad, kan vi säga, mellanfördomar och postjudice. Fördomar gör en bedömning innan du hartittat på fakta. Postjudice gör en bedömning i efterhand. Fördomär fruktansvärt, i den meningen att du begår orättvisor och du gör allvarmisstag. Postjudice är inte så hemskt. Du kan inte vara perfekt naturligtvis; dukan göra misstag också. Men det är tillåtet att göra en bedömning efter att duhar undersökt bevisen. I vissa kretsar är det även uppmuntras.
		-- Carl Sagan, The Burden of Skepticism, Skeptical Enquirer, Vol. 12, pg. 46

%
Om en person (a) är dåligt, (b) får behandling syftar till att göra honom bättre,och (c) blir bättre, då ingen kraft resonemang känt att den medicinska vetenskapen kanövertyga honom om att det inte kan ha varit den behandling som återställde hans hälsa.
		-- Sir Peter Medawar, The Art of the Soluble

%
Amerika har upptäckts tidigare, men det har alltid varit tystas ner.
		-- Oscar Wilde

%
Unix: Vissa säger att inlärningskurvan är brant, men du bara måste klättra det en gång.
		-- Karl Lehenbauer

%
Ibland, är för lång för lång.
		-- Joe Crowe

%
När dåliga män kombinera måste bra associera; annars kommer de att falla en efter en,en unpitied offer i en föraktlig kamp.
		-- Edmund Burke

%
Bakom allt den politiska retoriken som slungas mot oss från utlandet, vi äratt hämta hem en oantastlig faktum - [terrorism är] ett brott av alla civiliseradestandard, begåtts mot oskyldiga människor, bort från scenen av politiskakonflikt, och måste hanteras som ett brott. . . .   [I] n vår erkännande av arten av terrorism som ett brott ligger vår bästa hoppatt ta itu med det. . . .   [L] et oss använda de verktyg som vi har. Låt oss åberopa det samarbete vi harrätt att förvänta sig runt om i världen, och med detta samarbete låt oss krympade mörka och fuktiga områden av fristad tills dessa fega marodörer hållsatt svara som brottslingar i en öppen och offentlig rättegång för de brott de harbegåtts, och få det straff de så väl förtjänar.
		-- William H. Webster, Director, Federal Bureau of Investigation, 15 Oct 1985

%
"Av alla diktaturer som påverkar mänskligheten, är tyranni i religionen värst."
		-- Thomas Paine

%
"Jag säger att vi tar bort, nuke platsen från omlopp Det är det enda sättet att vara säker.."
		-- Corporal Hicks, in "Aliens"

%
"Det finns ingenting så dödligt som inte hålla upp till människor möjlighet attgör stora och underbara saker, om vi vill stimulera dem på ett aktivt sätt. "
		-- Dr. Harold Urey, Nobel Laureate in chemistry

%
"... Ordentlig uppmärksamhet till jordiska behoven hos de fattiga, den deprimerade ochförtryckta, naturligtvis skulle utvecklas från dynamisk, formulera, piggmedvetenhet om de stora målen för människor och samhälle han konspirerat för att resa. "
		-- David Baker, paraphrasing Harold Urey, in "The History of Manned Space Flight"

%
"Athens byggde Akropolis. Korinth var en handelsstad, är intresserade avrent materialistiska saker. Idag beundrar vi Aten, besöka den, bevaragamla tempel, men vi knappast någonsin satt sin fot i Korint. "
		-- Dr. Harold Urey, Nobel Laureate in chemistry

%
"Till stor del eftersom det är så konkret och spännande program och som sådan kommertjänar till att bevara intresset och entusiasmen hos hela spektrumet avsamhället ... Det är motiverad eftersom ... Programmet kan ge en känsla av gemensamtäventyr och prestation till samhället i stort. "
		-- Dr. Colin S. Pittendrigh, in "The History of Manned Space Flight"

%
Utmaningen för utforskning av rymden och i synnerhet av landnings män på månenrepresenterar den största utmaningen som någonsin har stått inför den mänskliga rasen. Ävenom det inte fanns några tydliga vetenskapliga eller andra argument för att fortsätta med dettauppgift, skulle hela historien om vår civilisation fortfarande förmå män mot denmål. Faktum är att monteringen av vetenskapliga och militären med dessa mänskligaargument skapar en så överväldigande fall att man kan bortse från endastdem som är blinda för de läror historia, eller som vill avbrytacivilisationens utveckling vid tidpunkten för största möjligheten och drama.
		-- Sir Bernard Lovell, 1962, in "The History of Manned Space Flight"

%
Idén om man lämnar denna jord och flyger till en annan himlakropp ochlandning där och kliva ut och gå över detta organ har en fascinationoch en drivande kraft som kan få landet till en nivå av energi, ambition,och kommer att jag inte ser i något annat företag. Jag tror att om vi ärärliga mot oss själva, måste vi erkänna att vi behövde att drivkraft extremtstarkt. Jag tror uppriktigt att rymdprogrammet, med sin bemannadelanda på månen, om klokt avrättades, blir spjutspets för enbred front av modiga och energiska aktiviteter på alla områdensträvan i det mänskliga sinnet - aktiviteter som inte kunde utförasutom i en mental klimat ambition och förtroende som sådan en spjutspetskan ge.
		-- Dr. Martin Schwarzschild, 1962, in "The History of Manned Space Flight"

%
Det mänskliga samhället - man i en grupp - reser sig ur sin dvala till nya nivåer avproduktiviteten endast under stimulans av djupt inspirerande och vanligenuppskattade mål. En slö världen tjänar ingen anledning väl; en pigg världarbetar hårt mot uppriktigt önskade mål ger möjlighet ochstyrkan mot vilken många ändar kan vara nöjd ... till oöverträffadsocial prestation.
		-- Dr. Lloyd V. Berkner, in "The History of Manned Space Flight"

%
Styrka i civiliserade samhällen bevaras av den utbredda känslan att högamål är lönande. Kraftfulla samhällen hyser en viss extravagansmål, så att män vandra förbi säkert tillhandahållande av personliggratifications. Alla starka intressen lätt bli opersonlig, kärleken bra väl utfört arbete. Det finns en känsla av harmoni om en sådan prestation,Peace väckts av något lönande.
		-- Alfred North Whitehead, 1963, in "The History of Manned Space Flight"

%
Jag tror inte att denna generation amerikaner är villig att avgå självatt gå till sängs varje kväll i ljuset av en kommunistisk måne ...
		-- Lyndon B. Johnson

%
Livet är densamma, med undantag för skor.
		-- The Cars

%
lila humBlandade bilarLaserljus, du tarAllt för att bevisaDu är på språngoch försvinnande
		-- The Cars

%
Kan vara du passerar den fina linjenEn dum förare slags ... off the wallDu håller den svalna när det är t-t täta... Ögonen öppna när du börjar falla.
		-- The Cars

%
Anpassa. Njut av. Överleva.
		-- The Cars

%
Fanns det färre dårar skulle knaves svälta.
		-- Anonymous

%
Mänskligheten har stjärnorna i sin framtid, och att framtiden är alltför viktigt att varaförlorade under bördan av ungdoms dårskap och okunnig vidskepelse.
		-- Isaac Asimov

%
Och publiken var stillas. En äldre man och undrade på den plötsliga tystnaden,vände sig till barn och bad honom att upprepa vad han hade sagt. Storögda,Barn höjde sin röst och sade återigen, "Varför har kejsaren ingenkläder! Han är naken! "
		-- "The Emperor's New Clothes"

%
"De som tror på astrologi lever i hus med grunderna förEnfaldigt Putty. "
		-- Dennis Rawlins, astronomer

%
Hittills har de definitiva slutsatser från Project Blue Book är:   1. ingen oidentifierat flygande föremål rapporteras, utreds och utvärderas      av flygvapnet någonsin gett någon indikation på hot mot vår      nationell säkerhet;   2. det har förekommit någon bevisning eller upptäcktes av Air      Kraft som siktats kategoriseras som OIDENTIFIERAD representerar      den tekniska utvecklingen eller principer utanför intervallet      dagens vetenskapliga rön; och   3. Det har inte funnits något bevis för att iakttagelser kategoriseras      som UNIDENTIFIED är utomjordiska fordon.- Sammanfattningen av Project Blue Book, en flygvapen studie av UFOn från 1950  till 1965, som citeras av James Randi i Flim-Flam!
		-- Dennis Rawlins, astronomer

%
De som tror att de tror på Gud, men utan passion i derashjärtan, utan ångest i åtanke, utan osäkerhet, utan tvekan,utan en del av förtvivlan även i deras tröst, tror endasti Gud idé, inte Gud själv.
		-- Miguel de Unamuno, Spanish philosopher and writer

%
Tvivel är en smärta för ensam för att veta att tro är hans tvillingbror.
		-- Kahlil Gibran

%
Tvivel är inte motsatsen till tro; Det är en del av tron.
		-- Paul Tillich, German theologian and historian

%
Tvivel är inte ett angenämt villkor, men säkerhet är absurd.
		-- Voltaire

%
Om bara Gud skulle ge mig några tydliga tecken! Som att göra en stor insättningi mitt namn på en schweizisk bank.
		-- Woody Allen

%
Jag kan inte bekräfta Gud om jag inte bekräfta man. Därför Jag försäkrar båda.Utan en tro på mänsklig enhet Jag är hungrig och ofullständig. mänsklig enhetär uppfyllelsen av mångfald. Det är harmoni av motsatser. Det ären många trängade struktur, med färg och djup.
		-- Norman Cousins

%
Att nedgradera det mänskliga sinnet är dålig teologi.
		-- C. K. Chesterton

%
... Meningsskiljaktigheter är advantageious i religion. De flera sekterutföra kontoret av en gemensam censor morum över varandra. är enhetlighetuppnåelig? Miljontals oskyldiga män, kvinnor och barn, sedankristendomens införande, har bränts, torterat, böter, fängelse;men vi har inte avancerat en tum mot enhetlighet.
		-- Thomas Jefferson, "Notes on Virginia"

%
Livet är en process, inte en princip ett mysterium levas, inte ett problem attlösas.
		-- Gerard Straub, television producer and author (stolen from Frank Herbert??)

%
Så vi följer våra irrande stigar och mycket mörkret fungerar som vår guide ochvåra tvivel tjänar till att lugna oss.
		-- Jean-Pierre de Caussade, eighteenth-century Jesuit priest

%
Tro kan definieras kortfattat som en ologisk tro på förekomsten avosannolik.
		-- H. L. Mencken

%
Och tror ni inte att ni alla kvinnor är en Eva? Guds dompå ditt kön uthärdar i dag; och med den alltid varar din positionkriminella i baren rättvisa.
		-- Tertullian, second-century Christian writer, misogynist

%
Jag bedöma en religion som bra eller dåligt beroende på om dess anhängarebli bättre människor som en följd av att öva det.
		-- Joe Mullally, computer salesman

%
Imitation är den ärligaste formen av plagiering.
		-- Joe Mullally, computer salesman

%
"Unibus timeout dödlig fälla programmet förlorade ledsen"
		-- An error message printed by DEC's RSTS operating system for the PDP-11

%
Hur många surrealist tar det att skruva i en glödlampa?En att hålla giraff och en för att fylla badkaret med färggladaelverktyg.
		-- An error message printed by DEC's RSTS operating system for the PDP-11

%
Hur många bayerska Illuminati tar det att skruva i en glödlampa?Tre: en att skruva fast den, och en att förvirra frågan.
		-- An error message printed by DEC's RSTS operating system for the PDP-11

%
Hur lång tid tar det en DEC servicetekniker att byta en glödlampa?Det beror på hur många dåliga han förde med sig.
		-- An error message printed by DEC's RSTS operating system for the PDP-11

%
Det gör mig någon skada för min granne att säga att det finns tjugo gudar eller ingen Gud.Det tar varken min ficka eller bryter benet.
		-- Thomas Jefferson

%
Jag tror inte på bekännelsen bekände av den judiska kyrkan, av den romerskaKyrka, av den grekiska kyrkan, av den turkiska kyrka, av den protestantiska kyrkan,eller av någon kyrka som jag känner till. Min egen uppfattning är min egen kyrka.
		-- Thomas Paine

%
Gud fordrar inte en enhetlighet i religion.
		-- Roger Williams

%
Den dagen kommer, då den mystiska generationen av Jesus, av Högsta väsendetsom Fadern, i livmodern av en jungfru kommer att klassificeras med fabeln omgenerering av Minerva i hjärnan hos Jupiter. Men vi får hoppas attgryning av förnuft och tankefrihet i dessa USA kommer att göra sig av meddenna artificiella ställningar och återställa till oss den primitiva och äktaläror detta mest vördade reformator av mänskliga misstag.
		-- Thomas Jefferson

%
Låt oss då medborgare, förena sig med ett hjärta och ett sinne. Låt ossåterställa till socialt umgänge som harmoni och kärlek utan vilkenfrihet och även livet självt är utan trista saker. Och låt oss reflekteraatt ha bannlyst från vårt land som religiös intolerans under vilkamänskligheten så länge blödde, har vi ännu fått lite om vi counternance enpolitisk intolerans som despotisk, som ond, och kan en bitter ochblodiga förföljelser.
		-- Thomas Jefferson

%
Jag finner inte i ortodox kristendom ett försonande drag.
		-- Thomas Jefferson

%
Jesu gudomlighet görs en bekväm täckmantel för absurditet. Ingenstans stans~~POS=HEADCOMPi evangelierna finner vi ett bud för bekännelser, bekännelsen, Eder,Lärdomar och hela carloads av andra dumt trumpery som vi finner iKristendom.
		-- John Adams

%
Bibeln är inte min bok och kristendom är inte min religion. jag skulle kunnaaldrig ge samtycke till de långa komplicerade rapporter Christian dogm.
		-- Abraham Lincoln

%
Som Jesus från Nasaret ... Jag tror att systemet med moral och hans religion,när han lämnade dem till oss, den bästa i världen någonsin sett eller sannolikt kommer att se;men jag uppfattar det har fått olika korrumperande ändringar och jag har,med de flesta av de nuvarande oliktänkande i England, några tvivel om hansgudomlighet.
		-- Benjamin Franklin

%
Jag skulle ha lovat de terrorister en resa till Disneyland om det skulle hablivit gisslan släppts. Jag tackar Gud att de var nöjda medmissiler och vi behövde inte gå till det extrema.
		-- Oliver North

%
Jag tror på en USA där separationen mellan kyrka och stat är absolut -där ingen katolsk prelat skulle berätta presidenten (han bör vara katolik)hur man ska agera, och ingen protestantisk präst skulle berätta för sina församlingsbor för vilkaatt rösta - där ingen kyrka eller kyrka skola beviljat några offentliga medel ellerpolitisk preferens - och där ingen människa nekas offentligt ämbete endasteftersom hans religion skiljer sig från president som kan utse honom ellermänniskor som kanske väljer honom.- Från John F. Kennedys tal till Greater Houston minister Association  September 12, 1960.
		-- Oliver North

%
Sanningen är att den kristna teologin, som alla andra teologi, är inte baramotsats till den vetenskapliga andan; det är också emot alla andra försökpå rationellt tänkande. Inte av en slump gör Genesis 3 gör faderkunskap en orm - slemmig, smyga och avskyvärda. Eftersom den tidigastedagar kyrkan som organisation har kastat sig våldsamt mot varjeförsök att befria kroppen och människans sinne. Det har varit, vid alla tidpunkter ochöverallt, vanliga och oförbätterlig försvarare av dåliga regeringar, dåliglagar, dåliga sociala teorier, dåliga institutioner. Det var under århundraden, enapologet för slaveri, eftersom det var apologet för den gudomliga nåde.
		-- H. L. Mencken

%
Uppfattningen att vetenskapen inte bryr sig om med första orsaker - att detlämnar fältet till teologi eller metafysik, och inskränker sig till enbarteffekter - detta begrepp har inget stöd i vanliga fakta. Om det kunde,vetenskap skulle förklara livets uppkomst på jorden på en gång - och det finnsall anledning att tro att det kommer att göra det på vissa inte alltför avlägsen i morgon.Att hävda att kunskapsluckor som möter sökaren måste fyllas,inte av patientens undersökning, utan genom intuition eller uppenbarelse, är helt enkelt att geokunnighet ett omotiverat och orimlig värdighet ....
		-- H. L. Mencken, 1930

%
Bevisen för känslor, utom i de fall då det har en stark målsättningstöd, är verkligen inga bevis alls, för varje igenkännbar känsla hardess motsats, och om man pekar ett sätt sedan en annan poäng åt andra hållet.Således känner argumentet att det finns en instinktiv längtan efter odödlighet,och att denna önskan visar sig vara ett faktum, blir puerile när det ärpåpekas att det finns också en kraftfull och utbredd rädsla för förintelse,och att denna fruktan, på samma princip visar att det inte finns någotbortom graven. Sådana barnsliga "bevis" är typiskt teologisk, ochde förblir teologiska även när de åberopas av män som gillar attsmickra sig genom att tro att de är vetenskapliga gents ....
		-- H. L. Mencken

%
Det finns i själva verket ingen anledning att tro att en viss naturfenomen,men underbart det kan tyckas i dag, kommer att finnas kvar för alltid oförklarligt.Förr eller senare de lagar som styr produktionen av livet självt kommer att varaupptäcktes i laboratoriet, och man kan etablera sig som en skapareför egen räkning. Saken verkligen är inte bara tänkbart; det äräven mycket sannolik.
		-- H. L. Mencken, 1930

%
Det bästa som vi kan göra är att vara vänlig och hjälpsam mot våra vänner ochmedpassagerare som klamrar sig fast på samma fläck av smuts medan vi ärdrivande sida vid sida för att vår gemensamma undergång.
		-- Clarence Darrow

%
Vi är här för att ge dig en dator, inte en religion.
		-- attributed to Bob Pariseau, at the introduction of the Amiga

%
... Kan det inte finnas någon offentlig eller privat stöd om grunden för åtgärden ärbruket av sanningen.
		-- George Jacob Holyoake

%
"Om ni ursäktar mig en minut, jag kommer att ha en kopp kaffe."- Sändning från Apollo 11: s LEM, "Eagle", till Johnson Space Center, Houston  20 juli 1969, 07:27
		-- George Jacob Holyoake

%
De ödmjuka bestrider viljan.
		-- George Jacob Holyoake

%
Jag är trött på att trampas på! Flädergudarna säger att de kan göra mig en man!Allt det kostar är min själ! Jag gör det, cuz nu är jag MAD !!!
		-- Necronomicomics #1, Jack Herman & Jeff Dee

%
   På Krat huvudskärm dök holo bilden av en man, och flera delfiner.Från mannens form, kunde Krat tala om det var en kvinna, troligen deras ledare.   "... Dumma varelser ovärdig namnet` sophonts. " Dåraktigt, pre-kännandeur sitt tvång; av vandrande mästare. Vi glida bort från alla dina väpnade styrka, skrattarpå din klumpighet! Vi glider bort som vi alltid kommer du patetiska varelser.Och nu när vi har en riktig försprång, kommer du aldrig fånga oss! vad bättrebevis för att stamceller gynnar inte dig, men oss! Finns det något bättre bevis ... "   Hån gick på. Krat lyssnade, rasande, men på samma gång savoringartisteri av det. Dessa män är bättre än jag trodde. deras förolämpningarär ordrik och uppblåst, men de har talang. De förtjänar heder, långsamdödsfall.
		-- David Brin, Startide Rising

%
"Jag är en genomsnittlig grön mor från yttre rymden"
		-- Audrey II, The Little Shop of Horrors

%
I likhet med mina föräldrar, jag har aldrig varit en vanlig församlingsmedlem eller churchgoer.Det verkar inte rimligt för mig att det är den typ av Gud somvakar över mänskliga angelägenheter, lyssnar till böner och försöker att styramänniskor att följa hans bud - det finns alldeles för mycket elände ochgrymhet för det. Å andra sidan, jag respekterar och avundas människorsom får inspiration från sina religioner.
		-- Benjamin Spock

%
Alla tillräckligt avancerad teknologi är omöjlig att skilja från en riggad demo.
		-- Andy Finkel, computer guy

%
Att vara schizofren är bättre än att leva ensam.
		-- Andy Finkel, computer guy

%
NowPrint. NowPrint. Clemclone, tillbaka till skuggorna igen.
		-- The Firesign Theater

%
Ja, många primitiva människor tror fortfarande denna myt ... Men i dagens teknisktvidden av framtiden, kan vi gissa som säkert saker var mycket annorlunda.
		-- The Firesign Theater

%
... Detta är en fantastisk syn. Hela rebell motstånd begravd under sexmiljoner inbundna exemplar av "The Naked Lunch".
		-- The Firesign Theater

%
Vi vill skapa dockor som drar sina egna strängar.
		-- Ann Marion

%
Jag vet ingenjörer. De älskar att förändra saker och ting.
		-- Dr. McCoy

%
På vår campus UNIX-systemet har visat sig vara inte bara en effektiv programvaraverktyg, men en agent för teknisk och social förändring inom universitetet.
		-- John Lions (University of New South Wales)

%
De som inte förstår Unix är dömda att uppfinna det, dåligt.
		-- Henry Spencer, University of Toronto Unix hack

%
"Du vet varför det finns så få sofistikerade terrorister i USAStaterna? Eftersom dina hackare har så mycket rörlighet i anläggningen.Här finns det ingen sådan rörlighet. Om du har det minsta intellektuellintegritet du inte kan stödja regeringen .... Det är därför den bästa datornsinnen tillhör oppositionen. "
		-- an anonymous member of the outlawed Polish trade union, Solidarity

%
"Varje Solidaritet centrum hade högar och högar av papper .... alla varäter papper och en polis var vid dörren. Allt du behöver göra är attböja en skiva. "- En anonym medlem av den förbjudna polska fackföreningen Solidaritet,  kommentera om fördelarna med att använda datorer för att stödja deras rörelse
		-- an anonymous member of the outlawed Polish trade union, Solidarity

%
Kläderna gör mannen. Nakna människor har liten eller ingen inverkan på samhället.
		-- Mark Twain

%
Ju tidigare alla djur är utdöda, desto snabbare kommer vi att hitta sina pengar.
		-- Ed Bluestone

%
Han är död, Jim.
		-- Ed Bluestone

%
New York ... när civilisationen faller sönder, minns vi var långt före dig.
		-- David Letterman

%
Du kan göra mer med ett vänligt ord och en pistol än med bara ett vänligt ord.
		-- Al Capone

%
Fontänen koden har skärpts något så att du inte längre kan doppa objekti en fontän eller dryck från en medan du svävar i luften på grund avlevitation.Teleportera till helvetet via en teleporte fälla kommer inte längre att uppstå omkaraktär inte har brandsäkerhet.
		-- README file from the NetHack game

%
Kom ihåg att det finns en stor skillnad mellan knä och böja.
		-- Frank Zappa

%
Jag tror att alla rättänkande människor i detta land är sjuka ochtrött på att höra att vanliga hyggliga människor är trötta på dettaland med att vara sjuk och trött. Jag är verkligen inte. Men jag ärtrött på att höra att jag är.
		-- Monty Python

%
"Det finns ingen preskriptionstid på dumhet."
		-- Randomly produced by a computer program called Markov3.

%
Det finns en tid i tidvatten män,Som var för vid översvämning, leder vidare till framgång.Å andra sidan, inte räkna med det.
		-- T. K. Lawson

%
För att följa dåraktiga prejudikat, och blinkningMed båda våra ögon, är lättare än att tänka.
		-- William Cowper

%
Det är kvalitet snarare än kvantitet som räknas.
		-- Lucius Annaeus Seneca (4 B.C. - A.D. 65)

%
Man kanske kan dividera om kvaliteten på ett enda experiment, ellerom sanningshalten i en viss försöks, men tar alla stödjandeexperiment tillsammans, är så stark sammanvägd lika lätt attförtjänar en klok man eftertanke.- Professor William Tiller, parapsychologist, Standford University,  kommentera psi forskning
		-- Lucius Annaeus Seneca (4 B.C. - A.D. 65)

%
Ingenting någonsin blir verklighet förrän den upplevs.
		-- John Keats

%
Din goda natur kommer att ge dig obegränsad lycka.
		-- John Keats

%
"Vår resa mot stjärnorna har utvecklats snabbt.1926 lanserade Robert Goddard första vätskegående raket,uppnå en höjd av 41 fot. 1962 John Glenn orbited jorden.1969, bara 66 år efter Orville Wright flög två fötter från marken12 sekunder, Neil Armstrong, Buzz Aldrin och jag höjden till måneni Apollo 11. "- Michael Collins   Tidigare astronaut och tidigare chef för National Air and Space Museum
		-- John Keats

%
De flesta människor uppvisar vad statsvetare kallar "konservatismbönderna. "Tappa inte vad du har. Ändra inte. Ta inte en chans,eftersom du kan hamna svälter ihjäl. Spela säkert. Köp lika mycketsom du behöver. Slösa inte tid.När vi tänker på risken, människor och företag inser i derashuvuden att riskerna är nödvändiga för att växa, för att överleva. Men när det kommer neratt hålla goda människor när kritan kommer, eller investera pengar inågot oprövad, bara de modiga nå djupt i sina fickor och spelaspelet som det måste spelas.
		-- David Lammers, "Yakitori", Electronic Engineering Times, January 18, 1988

%
"Vi kan inte schemalägga en orgie, det kan tolkas som slåss"
		-- Stanley Sutton

%
Helger gjordes för programmering.
		-- Karl Lehenbauer

%
"En gång hade han ett ben i Vita huset och nationen darrade under hansbrusar. Nu är han en SKRUTTIG påve i Coca-Cola bälte och en bror tillgivna pastorer som belabor halfwits i galvaniserat järn hyddor bakomjärnvägen varven. "- H.L. Mencken, skrivandet av William Jennings Bryan, ombud för supportrar  of Tennessee anti-evolution lag på omfattningar "Monkey Trial" i 1925.
		-- Karl Lehenbauer

%
... Vi måste motsats den överväldigande dom från konsekventobservationer och slutsatser i tusental. Jorden är miljarderår gammal och dess levande varelser är förenade genom band av evolutionärahärkomst. Forskare anklagas för att främja dogmer genom så anger, mengör vi helt folk intolerant när de förkunnar att jorden är varkenflata eller i mitten av universum? Vetenskap * har * lärt oss någrasaker med tillförsikt! Evolution på en forntida jord är ocksåetablerades som vår planets form och position. Vår fortsatta kampatt förstå hur evolutionen händer (det "evolutionsteorin") intekasta vår dokumentation av dess förekomst - den "faktum evolution" -sättas.- Stephen Jay Gould, "The Bedömning på kreationism", The Skeptical Inquirer,  Vol XII No. 2
		-- Karl Lehenbauer

%
Detta var den ultimata formen av flärd bland teknik freaks - att haett system så komplett och sofistikerade att ingenting visade; inga maskiner,inga sladdar, inga kontroller.
		-- Michael Swanwick, "Vacuum Flowers"

%
Män borde veta att endast från hjärnan och från hjärnan uppstår vårnöjen, glädje, skratt och skämt samt våra sorger, smärtor, sorgeroch tårar. ... Det är samma sak som gör oss galna eller yrande, inspireraross med fruktan och rädsla, antingen genom natt eller dag, ger oss sömnlöshet,olämpliga misstag, planlösa oro, tankspriddhet och handlingar som äri strid med vana ...
		-- Hippocrates (c. 460-c. 377 B.C.), The Sacred Disease

%
Modern psykologi tar helt för givet att beteende och neural funktionär perfekt korrelerade, är att en helt orsakad av den andra. Det finnsingen separat själ eller livskraft att hålla ett finger i hjärnan då och då ochgör neurala celler gör vad de annars inte skulle. Faktiskt, naturligtvis, dettaär bara en arbetshypotes .... Det är fullt tänkbart att en dag iantagande måste avvisas. Men det är också viktigt att se till att vihar inte nått den dagen ännu: arbetshypotesen är en nödvändig en ochDet finns inga riktiga bevis motsätter sig det. Vårt misslyckande att lösa ett problem sålångt inte gör det olösligt. Man kan inte logiskt vara en deterministisk ifysik och biologi, och en mystisk i psykologi.
		-- D. O. Hebb, Organization of Behavior:  A Neuropsychological Theory, 1949

%
Förhärskande tro att kunskap kan utnyttjas från tidigare inkarnationer ellerfrån en "universell sinne" (förvaret av alla tidigare visdom och kreativitet)inte bara är osannolikt men också orättvist förnedra den fantastiska prestationerindividuella mänskliga hjärnor.- Barry L. Beyerstein, "Hjärnan och medvetande: Inblandning för Psi  Fenomen ", The Skeptical Inquirer, Vol. XII nr 2, PPG. 163-171
		-- D. O. Hebb, Organization of Behavior:  A Neuropsychological Theory, 1949

%
... Lyckligtvis är ansvaret för att tillhandahålla bevis på den del avden person som gör anspråk, inte kritikern. Det är inte ansvaretUFO skeptiker att bevisa att ett UFO aldrig har funnits, inte heller är detansvar paranormala-hälsa-skade skeptiker att bevisa att kristallereller färgade ljus läkt aldrig någon. Skeptiker roll är att påpekapåståenden som inte är tillräckligt stöds av godtagbara bevis ochtillhandahålla rimliga alternativa förklaringar som är mer i linje medden accepterade vetenskapliga bevis. ...
		-- Thomas L. Creed, The Skeptical Inquirer, Vol. XII No. 2, pg. 215

%
"Ada är ett verk av en arkitekt, inte datavetare."
		-- Jean Icbiah, inventor of Ada, weenie

%
Otroliga påståenden kräver extraordinära bevis. Det finns många exempel påutomstående som så småningom störtade inrotade vetenskapliga ortodoxier, mende segrade med obestridliga data. Oftare flagranta rön sommotsäger väletablerad forskning visar sig vara artefakter. jag harhävdade att acceptera psykiska krafter, reinkarnation, "kosmiskt medvetande"och liknande, skulle innebära grundläggande ändringar av grunderna förneurovetenskapen. Innan överge materialistiska teorier om sinnet som har betalatvacker utdelning, bör vi insistera på bättre bevis för psi fenomenän finns närvarande, särskilt när neurologi och psykologi självaerbjuda mer trovärdiga alternativ.- Barry L. Beyerstein, "Hjärnan och medvetande: Inblandning för Psi   Fenomen ", The Skeptical Inquirer, Vol. XII nr 2, PPG. 163-171
		-- Jean Icbiah, inventor of Ada, weenie

%
Evolution är en bankrutt spekulativ filosofi, inte ett vetenskapligt faktum.Endast en andligt konkurs samhälle någonsin kunde tro det. ... Endastateister kan acceptera detta Satanic teori.
		-- Rev. Jimmy Swaggart, "The Pre-Adamic Creation and Evolution"

%
Evolution är lika mycket ett faktum som jorden slå på sin axel och går runtsolen. Vid ett tillfälle detta kallades Kopernikus teori; men närbevis för en teori blir så överväldigande att ingen informerade personenkan tvivlar på det, är det brukligt för forskare att kalla det ett faktum. Att allanuvarande liv härstammar från tidigare former, över stora sträckor av geologiskatid, är så fast etablerad som Copernican kosmologi. biologer skiljerendast med avseende på teorier om hur processen fungerar.- Martin Gardner, "Irving Kristol och fakta av liv",   Den Skeptical Inquirer, Vol. XII No. 2, ppg. 128-131
		-- Rev. Jimmy Swaggart, "The Pre-Adamic Creation and Evolution"

%
... Det är tråkigt att hitta honom belaboring vetenskapssamhället för sin enademotstånd mot okunniga kreation som vill lärare och läroböcker tillge lika mycket tid att skruva argument som har framförts inte ett steg längreden Flyblown retorik biskop Wilberforce och William Jennings Bryan.- Martin Gardner, "Irving Kristol och fakta av liv",   Den Skeptical Inquirer, Vol. XII No. 2, ppg. 128-131
		-- Rev. Jimmy Swaggart, "The Pre-Adamic Creation and Evolution"

%
... Boken är värd uppmärksamhet för bara två skäl: (1) den angriperförsök att avslöja falska paranormala studier; och (2) det är mycket bra ochrimligen skrivit och så snarare svårare att avfärda eller vederlägga genom enkelhånfull.- Harry Eagar, granska "Beyond the Quantum" av Michael Talbot,   Den Skeptical Inquirer, Vol. XII No. 2, ppg. 200-201
		-- Rev. Jimmy Swaggart, "The Pre-Adamic Creation and Evolution"

%
Nu lägger jag mig ner för att sovaJag hör sirenerna på gatanAlla mina drömmar är gjorda av kromJag har inget sätt att få tillbaka hem
		-- Tom Waits

%
Jag är här med folkviljan och jag kommer inte att lämna tills jag får min regnrocktillbaka.
		-- a slogan of the anarchists in Richard Kadrey's "Metrophage"

%
Hur många kärnkraftsingenjörer tar det att byta en glödlampa?Sju: En för att installera den nya glödlampan, och sex för att bestämma vad man ska göra        med den gamla en för de kommande 10.000 år.
		-- a slogan of the anarchists in Richard Kadrey's "Metrophage"

%
Mike lag:För en timmer företag som sysselsätter två män och en cut-off såg, demarginalprodukt av arbetskraft för ett obegränsat antal ytterligare arbetskraftär lika med noll tills förvärvet av en annan cut-off såg.Låt oss inte ens överväga en motorsåg.- Mike Dennison[Du kan alltid schema sågen, men - red.]
		-- a slogan of the anarchists in Richard Kadrey's "Metrophage"

%
Så länge vi kommer att uppfinna hjulet igen, kan vi lika gärna försöka göradet runda denna gång.
		-- Mike Dennison

%
Denna kombination av en enorm militära etablissemanget och en stor armarindustrin är nu i den amerikanska erfarenheten ... Vi får inte misslyckas med attförstå dess allvarliga konsekvenser ... Vi måste skydda sig motförvärv av obefogad påverkan ... av militär-industriellakomplex. Potentialen för den katastrofala ökningen av missriktad kraftexisterar och kommer att bestå.
		-- Dwight D. Eisenhower, from his farewell address in 1961

%
Denna restaurang var reklam frukost helst. Så jag beställdefrench toast i renässansen.
		-- Steven Wright, comedian

%
Alla har en mening med livet. Kanske din är att titta på tv.
		-- David Letterman

%
En hel del av de saker jag gör är så minimal, och det är utformat för att vara minimal.Komponenten det är vad som är attraktivt. Det är konstigt, för det är såintellektuellt lamt. Det är svårt att se mig göra det för resten avmitt liv. Men samtidigt är det vad jag gör bäst.
		-- Chris Elliot, writer and performer on "Late Night with David Letterman"

%
e-trovärdighet: icke-guaranteeable sannolikheten för att elektroniskt datadu ser är äkta snarare än någon är påhittade skit.
		-- Karl Lehenbauer

%
När folk är överens med mig, jag tror alltid att jag måste vara fel.
		-- Oscar Wilde

%
Min mamma är en fisk.
		-- William Faulkner

%
Ju längre den andliga utvecklingen av mänskligheten framsteg, desto mer säker på att dettycks mig att vägen till äkta religiositet inte ligger genomrädsla för livet, och rädslan för döden, och blind tro, utan genom att strävaefter rationell kunskap.
		-- Albert Einstein

%
Ju mer en människa präglas av beställda korrekthet alla händelser, desto fastareblir hans övertygelse om att det inte finns något utrymme kvar vid sidan av detta beordraderegelbundenhet för orsakerna till en annan karaktär. För honom varken regeln ommänsklig eller regeln om gudomliga viljan existerar som en oberoende orsak till naturlighändelser. För att vara säker, läran om en personlig Gud störa naturligahändelser kan aldrig vederläggas, i egentlig mening, av vetenskapen, för dettadoktrin kan alltid ta sin tillflykt i de områden där vetenskaplig kunskaphar ännu inte kunnat sätta sin fot.Men jag är övertygad om att ett sådant beteende på den del av företrädarnareligionens skulle inte bara vara ovärdig men också dödlig. För en doktrin somkan bibehålla sig inte klart ljus, men endast i mörker, kommerav nödvändighet förlorar sin effekt på mänskligheten, med oöverskådliga skador på människorsframsteg. I sin kamp för etisk bra, religionsläraremåste ha resning att ge upp läran om en personlig Gud, det vill sägage upp den källa till rädsla och hopp som tidigare placerade så stortbefogenheter i händerna på prästerna. I sitt arbete som de kommer att behöva utnyttjasig av de krafter som kan odla det goda, detDet är sant, och det sköna i mänskligheten själv. Detta är, för att vara säker, en mersvårt men en ojämförligt mer värdig uppgift.
		-- Albert Einstein

%
Någon som vet historia, särskilt Europas historia, kommer, tror jag,inse att dominansen av utbildning eller regerings av någonsärskild religiös tro är aldrig en glad arrangemang för människor.
		-- Eleanor Roosevelt

%
De flesta icke-katoliker vet att katolska skolor gör en störreservice till vår nation än de offentliga skolor där omstörtande läroböckerhar använts, i vilken kommunist sinnade lärare har undervisat, och frånvars klassrum Kristus och även Gud själv är spärrade.
		-- from "Our Sunday Visitor", an American-Catholic newspaper, 1949

%
De av oss som tror på rätten för varje människa att tillhöra vadkyrka han anser det lämpligt, och att dyrka Gud på sitt eget sätt, kan inte klandrasfördomar när vi inte vill se statlig utbildning i samband medreligiösa kontroll av skolor, som betalas av skattebetalarnas pengar.
		-- Eleanor Roosevelt

%
Andligt ledarskap bör förbli andligt ledarskap och tidsmakt bör inte bli alltför viktig i någon kyrka.
		-- Eleanor Roosevelt

%
Sanningen har alltid visat sig främja bästa för mänskligheten ...
		-- Percy Bysshe Shelley

%
Om ateism är att användas för att uttrycka sinnesstämning i vilken Gud äridentifierad med unknowable, och teologi uttalas att vara ensamling av meningslösa ord om obegripliga chimärer, sedanJag har inga tvivel om, och jag tror att få människor tvivlar, att ateister ärrikligt som björnbär ...
		-- Leslie Stephen (1832-1904), literary essayist, author

%
Det är fel alltid, överallt och för alla att tro något påtillräckliga bevis.
		-- W. K. Clifford, British philosopher, circa 1876

%
Varför, när ingen ärlig man kan förneka privat att varje ultimata problemet ärinsvept i den djupaste mysterium, gör ärliga män förkunna i predikstolarsom tveklöst säkerhet åligger de mest dåraktiga och okunniga?Är det inte ett spektakel att änglarna skratta? Vi är ett företag medokunniga varelser, känner oss igenom dimma och mörker, bara lärandevara oupphörligt upprepas misstag, få en glimt av sanningenfalla in alla tänkbara fel, svagt kräsna tillräckligt lätt förvåra dagliga behov, men hopplöst skiljer sig när vi försöker att beskrivaden ultimata ursprung eller slutet av våra vägar; Och ändå, när en av oss venturesatt förklara att vi inte vet karta över universum liksom kartanav vår oändligt socken, han tutade, avskydda och kanske höra atthan kommer bli fördömd i all evighet för hans trolöshet ...
		-- Leslie Stephen, "An agnostic's Apology", Fortnightly Review, 1876

%
Tills dess får vi nöja oss med att erkänna öppet, vad du (religionists)viska i din andedräkt eller gömma sig i teknisk jargong, att den gamlaHemligheten är en hemlighet fortfarande; att man vet ingenting om det oändliga ochAbsolut; och att veta någonting, han hade bättre att inte vara dogmatisk omhans okunnighet. Och under tiden kommer vi att sträva efter att vara så välgörande sommöjligt, och medan du trumpet fram officiellt din förakt för vårskepsis, kommer vi åtminstone försöka att tro att du åläggsav din egen rasa.
		-- Leslie Stephen, "An agnostic's Apology", Fortnightly Review, 1876

%
Förbindelse är den enda äventyr öppna för feg.
		-- Voltaire

%
Vad är tolerans? - Det är en följd av mänskligheten. Vi är alla bildadeav svaghet och fel; Låt oss förlåta ömsesidigt varandras dårskap -det är det första naturens lag.
		-- Voltaire

%
Det är uppenbart att den person som förföljer en man, hans bror, eftersomhan är inte av samma åsikt, är ett monster.
		-- Voltaire

%
Jag försöker bara att hjälpa till att låta ljuset av historiska sanningen i detruttnande massa utsliten tanke som fäster den moderna världenmedeltida föreställningar om kristendomen och som lever fortfarande bland oss ​​-en allvarligaste hindret för religion och moral, och ett hot mot helanormal utveckling av samhället.
		-- Andrew D. White, author, first president of Cornell University, 1896

%
Mannen knappa liv som inte är mer godtrogen än han borde vara .... Detnaturlig disposition är alltid att tro. Det förvärvas visdom och erfarenhetbara att lära misstro, och de mycket sällan lär det nog.
		-- Adam Smith

%
Jag satte hagelgevär i en Adidas väska och vadderad ut med fyra par tennisstrumpor, inte min stil alls, men det var vad jag siktar på: Om de trordu är rå, gå tekniskt; om de tror att du är tekniskt, gå rå. Jag är enmycket teknisk pojke. Så jag bestämde mig för att få så rå som möjligt. Dessa dagar,Men du måste vara ganska teknisk innan du ens kan aspirera påråhet.
		-- Johnny Mnemonic, by William Gibson

%
Men på religiösa frågor kan det vara liten eller ingen kompromiss.Det finns ingen plats där människor är så fast som deras religiösaövertygelser. Det finns ingen mer kraftfull allierad en kan göra anspråk på en debatt änJesus Kristus, eller Gud, eller Allah, eller vad man kallar det högsta väsen.Men precis som alla kraftfulla vapen, användningen av Guds namn på en räkningbör användas sparsamt. De religiösa fraktioner som växerhela vårt land inte använder sin religiösa inflytande med visdom.De försöker tvinga statsledningen till efter deras ställning100 procent. Om du inte håller med dessa religiösa grupper på ettsärskilt moralisk fråga, de klagar, de hotar dig med en förlust avpengar eller röster eller båda. Jag är uppriktigt trött på den politiskapredikanter över detta land talar om för mig som medborgare att om jag vill varaen moralisk person, måste jag tro på "A", "B", "C" och "D" Precis som görde tror att de är? Och varifrån har de antar att göra anspråk pårätt att diktera sina moraliska övertygelser för mig? Och jag är ännu mer arg somen lagstiftare som måste utstå hot om varje religiös grupp somtror att det har någon Gud beviljas rätten att kontrollera min röst på varje rullering i senaten. Jag varnar dem idag: Jag kommer att kämpa dem allasteg på vägen om de försöker att diktera sina moraliska övertygelser för allaAmerikaner i namn av "konservatism".
		-- Senator Barry Goldwater, from the Congressional Record, September 16, 1981

%
"Jag tror att varje god kristen borde sparka Falwell ass."- Senator Barry Goldwater, på frågan vad han tyckte om Jerry Falwell: sförslag om att alla goda kristna bör vara mot Sandra Day O'Connornominering till Högsta domstolen
		-- Senator Barry Goldwater, from the Congressional Record, September 16, 1981

%
... Och ingen filosofi, tyvärr har alla svaren. Oavsett hur säkervi kan vara om vissa aspekter av vår tro, det finns alltid smärtinkonsekvenser, undantag och motsägelser. Detta är sant i religionen somdet är i politik, och är självklart att alla utom fanatiker och den naiva.När det gäller fanatiker, vars antal är legio i vår egen tid, kanske vi vararekommenderas att lämna dem till himlen. De kommer inte, tyvärr, gör osssamma artighet. De attackerar oss och varandra, och oavsettprotester till fredliga avsikter, gör blodiga rekord av historien klaratt de lätt är anordnade för att återställa till svärdet. Min egen tro påGud, då är just det - en fråga om tro, inte kunskap. Min respektför Jesus Kristus härrör från det faktum att han tycks ha varitmest dygdiga invånare i planeten jorden. Men även välutbildade kristnaär frustrerade i sin törst efter visshet om den älskade figurJesus på grund av den obestridliga tvetydigheten i bibliska rekord.En sådan tvetydighet är inte uppenbart för barn eller fanatiker, men varjeerkända bibelkännare är fullt medveten om det. En del kristna, tyvärr,gripa formell liggande för att dölja en sådan verklighet.- Steve Allen, komiker, från en essä i boken "mod  Övertygelse ", redigerad av Philip Berman
		-- Senator Barry Goldwater, from the Congressional Record, September 16, 1981

%
... Det är fortfarande sant att en uppsättning av kognitiva föreställningar omGuds existens i någon igenkännbar mening kontinuerlig med den storasystem i det förflutna, religiösa läror utgör en spekulativhypotesen om en extremt låg ordning av sannolikhet.
		-- Sidney Hook

%
En fanatiker är en person som inte kan ändra sig och kommer inte att byta ämne.
		-- Winston Churchill

%
Vi kämpar mot humanism, vi kämpar mot liberalismen ...vi kämpar mot alla system av Satan som förstörvår nation idag ... vår kamp är med Satan själv.
		-- Jerry Falwell

%
De [predikanter] fruktar före vetenskapen som häxor gör tillvägagångssättetdagsljus och bister uppsyn på den ödesdigra förebud tillkännage subversionsav duperies där de bor.
		-- Thomas Jefferson

%
Heliga bör alltid bedömas skyldig tills de bevisats oskyldiga.
		-- George Orwell

%
Som jag argumenterade i "älskade Son", en bok om min son Brian och motivetreligiösa kommuner och kulter, ett resultat av korrekt tidig instruktioni förfarandena enligt rationellt tänkande kommer att vara att göra plötsliga meningslösaomvandlingar - till någonting - mindre troligt. Brian inser nu detta ochhar efter elva år, lämnade sekt han var förknippad med. DeProblemet är att när ett otränat sinne har gjort ett formellt åtagande atten religiös filosofi - och det spelar ingen roll om den filosofinär i allmänhet rimliga och hög sinnade eller fullständigt bisarra ochirrationella - befogenheter anledning är förvånansvärt ineffektiva iförändra den troendes sinne.- Steve Allen, komiker, från en essä i boken "mod  Övertygelse ", redigerad av Philip Berman
		-- George Orwell

%
Ingenting är lättare än att fördöma missdådaren; ingenting är svårareän att förstå honom.
		-- Fyodor Dostoevski

%
Vi kanske inte kan övertyga hinduer att Jesus och inte Vishnu börstyra sin andliga horisont, eller muslimer som Buddha är påcentrum för deras andliga universum, eller hebréer att Muhammed är en storprofet, inte heller de kristna som Shinto bäst uttrycker sin andligaoro, för att inte tala om det faktum att vi inte kan fåKristna att komma överens sinsemellan om deras förhållande till Gud.Men alla kommer att enas om ett förslag som de har djup andligresurser. Om dessutom kan vi få dem att acceptera ytterligarepåståendet att oavsett vilken form Gudomen kan ha sin egen teologi,Gudomen är inte bara yttre, men inre och verkar genom dem, ochde själva ge bevis eller vederlägga Gudomen i vad de gör ochtror; om denna ytterligare förslag kan godtas, då kommer vi attmycket närmare till en verkligt religiösa situationen på jorden.
		-- Norman Cousins, from his book "Human Options"

%
Messias kommer. Det kommer att finnas en uppståndelse från de döda - allade saker som judarna trodde på innan de fick så jävla sofistikerad.
		-- Rabbi Meir Kahane

%
Världen är ingen plantskola.
		-- Sigmund Freud

%
Om man frågar varför den amerikanska traditionen är så stark mot allaanslutning av kyrka och stat, varför det fruktar även grunderna ireligionsundervisning i statliga underhållna skolor, omedelbar ochytliga svar är inte långt att söka ....Orsaken låg i stort sett i mångfald och vitalitet av de olikavalörer, varje ganska säker på att, med en rättvis fält och ingen fördel,det kan göra sin egen väg; och varje animerad av en svartsjuk rädsla för att,Om någon anslutning av stat och kyrka tilläts vissa rivalvalör skulle få en otillbörlig fördel.- John Dewey (1859-1953), amerikansk filosof,  från "Demokrati i skolorna", 1908
		-- Sigmund Freud

%
Redan andan i vår skolgång genomsyras med en känsla av attvarje ämne, varje ämne, varje själva verket måste varje professed sanning varagenomgå en viss publicitet och opartiskhet. alla erbjudnaprover av lärande måste gå till samma analys-rum och utsättas förgemensamma tester. Det är kärnan i alla dogmatiska religioner att anse atten sådan "show-down" är vanhelgande och pervers. det karakteristiskareligion, från deras synvinkel, är att det är intellektuellthemlighet, inte offentliga; egendomligt avslöjat, i allmänhet inte känt;auktoritativt förklarade inte kommuniceras och testas i vanligasätt ... Det är relevant att påpeka att så länge som religion ärtänkt som det är nu av den stora majoriteten av bekännande religionists,finns det något motsägelsefullt att tala om utbildning ireligion i samma mening som vi talar om utbildning i ämnendär metoden för fri utredning har gjort sin väg. "Religiösa"skulle vara den sista att vara beredd att antingen historiainnehållet i religion bör läras ut i denna anda; medan detill vilken vetenskaplig synpunkt är inte enbart en teknisk anordning,men är förkroppsligandet av integritet åtanke måste protestera motdess undervisas i någon annan anda.- John Dewey (1859-1953), amerikansk filosof,  från "Demokrati i skolorna", 1908
		-- Sigmund Freud

%
I den breda och sista mening alla institutioner är pedagogiska imeningen att de arbetar för att bilda attityder, dispositioner, förmågoroch funktionshinder som utgör en konkret personlighet ... om dettauppfostrande processen bedrivs i en övervägande demokratisk eller ickedemokratiskt sätt blir därför en fråga om transcendent betydelseinte bara för själva utbildningen men för dess slutliga effekt på allaintressen och aktiviteter i ett samhälle som har åtagit sig att den demokratiskalivsstil.
		-- John Dewey (1859-1953), American philosopher

%
Historien visar att det mänskliga sinnet, matas med konstant anslutningarna av kunskap,periodvis blir för stor för sin teoretiska beläggningar, och bristerdem sönder visas i nya habiliments, som utfodring och växandegrub, med jämna mellanrum, kastar sin alltför snäv hud och förutsätter en annan ...Verkligen imago människans tillstånd verkar vara oerhört avlägsen, men varjeruggning är ett steg som gjorts.
		-- Charles Darwin, from "Origin of the Species"

%
... Jag skulle vilja gå så långt som att föreslå att, om det inte vore för vårt ego ochsträvan att vara annorlunda, skulle de afrikanska apor ingå i vårfamilj, Hominidae.
		-- Richard Leakey

%
Det är otänkbart att en omdömesgill observatör från ett annat solsystemskulle se i vår art - som har tenderat att vara grym, destruktiva,slösaktig och irrationella - kronan och toppen av kosmiska evolutionen.Tittar oss som kulmen på * något * är grotesk; visning osssom en övergångs art är mer förnuftigt - och ger oss mer hopp.- Betty McCollister, "Våra Övergångs Species",  Fritt få undersöka magazine, Vol. 8, nr 1
		-- Richard Leakey

%
"Jo, du ser, det är en övergångs varelse. Det är en pissa fattigareptil och inte så mycket av en fågel. "- Melvin Konner, från "Tangled Wing", citerar en zoolog som harstuderade archeopteryx och fann det "mycket som människor"
		-- Richard Leakey

%
"Du behöver kärleksfull omsorg en gång i veckan - så att jag kan smälla dig i form."
		-- Ellyn Mustard

%
"Det kan vara så att vår roll på denna planet är inte att dyrka Gud utan skapa honom. "
		-- Arthur C. Clarke

%
"Varför ska vi subventionera intellektuell nyfikenhet?"
		-- Ronald Reagan

%
"Det finns inget nytt under solen, men det finns massor av gamla saker Vi vet inte ännu. "
		-- Ambrose Bierce

%
"Plan för att kasta en bort. Du kommer i alla fall."
		-- Fred Brooks, "The Mythical Man Month"

%
Du behöver kärleksfull omsorg en gång i veckan - så att jag kan smälla dig i form.
		-- Ellyn Mustard

%
"Det kan vara så att vår roll på denna planet är inte att dyrka Gud utan skapa honom. "
		-- Arthur C. Clarke

%
"Varför ska vi subventionera intellektuell nyfikenhet?"
		-- Ronald Reagan

%
"Det finns inget nytt under solen, men det finns massor av gamla saker Vi vet inte ännu. "
		-- Ambrose Bierce

%
Mellanöstern är förvisso kopplingen av oron för en lång tid framöver -med skiftande aktörer, men samma spel: omvälvning. Jag tror att vi kommer att varakonfrontera militant islam - särskilt nedfall från den iranskarevolution - och religion kommer ännu en gång, eftersom det har i vår egen meravlägsna förflutna - spela en roll åtminstone som fanbärare i död och förödelse.- Bobby R. Inman, amiral, USN, Pensionerad, tidigare chef för Naval Intelligence,  vice chef för DIA, tidigare chef för NSA, biträdande chef för  Central Intelligence, tidigare ordförande och VD för MCC.
		-- Ambrose Bierce

%
... En sak är att, till skillnad från alla andra västerländska demokrati som jag känner till,detta land har fungerat sedan dess början med en grundläggande misstroregering. Vi utgörs inte för effektiv drift av regeringen,men för att minimera risken för maktmissbruk. Det tog händelsernaav Roosevelt eran - en katastrofal ekonomisk kollaps och ett världskrig -att införa den starka staten som vi nu vet. Men i de flestadelar av landet i dag, är motvilja mot att ha regeringen fortfarandestark. Jag tror, ​​spärra en rad katastrofala händelser, som vi kanse till åtminstone ett decennium under vilket många av de stora problemenrunt detta land måste behandlas på annat sätt än institutionerfederala regeringen.- Bobby R. Inman, amiral, USN, Pensionerad, tidigare chef för Naval Intelligence,  vice chef för DIA, tidigare chef för NSA, vice katalog  Central Intelligence, tidigare ordförande och VD för MCC.[De statist yttranden här är inte de kakan redaktör -ED.]
		-- Ambrose Bierce

%
"Jag har bara ett ord för dig, min pojke ... plast."
		-- from "The Graduate"

%
"Det finns en sådan fin linje mellan geni och dumhet."
		-- David St. Hubbins, "Spinal Tap"

%
"Om Diet Coke inte fanns skulle det ha varit nödvändigt att uppfinna den."
		-- Karl Lehenbauer

%
Jag närmade sig med de motsatta synpunkter och råd, och av män somär lika säker på att de representerar den gudomliga viljan. Jag är säker på attantingen det ena eller det andra är fel i tron, och kanske i vissaavseenden, båda.Jag hoppas att det inte kommer att vara vanvördig av mig att säga att om det är sannolikt attGud skulle avslöja sin vilja till andra på en punkt så förbunden med min plikt,det kan antas att han skulle avslöja det direkt till mig.
		-- Abraham Lincoln

%
I rymden kan ingen höra dig fisa.
		-- Abraham Lincoln

%
Hjärnskador är allt i huvudet.
		-- Karl Lehenbauer

%
Önskar och hoppas lyckas kräsna tecken på naturlighet där förnuft ochnoggrann vetenskapligt förfarande misslyckas.
		-- James E. Alcock, The Skeptical Inquirer, Vol. 12

%
"Det är bättre att ha försökt och misslyckats än att ha misslyckats med att prova, menResultatet är detsamma. "
		-- Mike Dennison

%
"Skapande vetenskap" har inte skrivit läroplanen av en anledning så enkeloch så grundläggande att vi ofta glömmer att nämna det: eftersom det är falskt, ocheftersom goda lärare förstå exakt varför det är falskt. Vad kan varamer destruktivt av det mest ömtåliga men mest värdefull resurs i vårHela intellektuella arv - god undervisning - än ett lagförslag som tvingarärade lärare att smutsa deras heliga förtroende genom att ge lika behandlingtill en doktrin inte bara kända för att vara falsk, men beräknas att underminera någonallmän förståelse för vetenskap som ett företag?
		-- Stephen Jay Gould, "The Skeptical Inquirer", Vol. 12, page 186

%
Det är inte bra att ses som en som ödmjukt underkastar sig fräckhet ochskrämsel.
		-- Stephen Jay Gould, "The Skeptical Inquirer", Vol. 12, page 186

%
"Oberoende av gällande hastighetsgräns, din Buick måste drivas påhastigheter snabbare än 85 MPH (140kph). "
		-- 1987 Buick Grand National owners manual.

%
"Din attityd avgör din inställning."
		-- Zig Ziglar, self-improvement doofus

%
Att argumentera att de nuvarande teorier om hjärnans funktion misstänkliggöra ESP,Telekinesi, reinkarnation, och så vidare, jag ofta utmanas medden mest populära av alla neuro mytologier - den uppfattningen att vi normaltAnvänd endast 10 procent av våra hjärnor ...Denna "cerebral reservdäck" -konceptet fortsätter att ge näring åt kundkrets"pop psykologer" och deras många system självförbättring återvinning. Somen metafor för det faktum att några av oss till fullo utnyttja våra talanger, som kundeförneka det? Som en fristad för ockultister som söker ett neuralt grund av den mirakulösa,det lämnar mycket övrigt att önska.- Barry L. Beyerstein, "Hjärnan och medvetande: Inblandning för   Psi Phenomena ", The Skeptical Enquirer, Vol. XII, nr 2, sid. 171
		-- Zig Ziglar, self-improvement doofus

%
Thufir är en Harkonnen nu.
		-- Zig Ziglar, self-improvement doofus

%
"Genom lång tradition, jag tar tillfället i akt stund andradesigners i tunn förklädnad av god, ren kul. "
		-- P. J. Plauger, from his April Fool's column in April 88's "Computer Language"

%
"Om du vill äta flodhäst, you got att betala frakten."
		-- attributed to an IBM guy, about why IBM software uses so much memory

%
Parkinsons lag: Arbete expanderar för att fylla tiden anvisade det.
		-- attributed to an IBM guy, about why IBM software uses so much memory

%
Karls version av Parkinsons lag: Arbete expanderar överskrida tiden anvisade det.
		-- attributed to an IBM guy, about why IBM software uses so much memory

%
Det är bättre att aldrig har provat något än att ha provat något ochmisslyckades.
		-- motto of jerks, weenies and losers everywhere

%
"Våra resor till stjärnorna kommer att göras på rymdskepp som skapats av beslutsamma,hårt vetenskapsmän och ingenjörer som tillämpar principerna om vetenskap, inteombord flygande tefat styrda av små grå utomjordingar från en annan dimension. "- Robert A. Baker, "The Aliens bland oss: hypnotisk regression Revisited",   Den Skeptical Inquirer, Vol. XII, nr 2
		-- motto of jerks, weenies and losers everywhere

%
"... Alla goda data mönster bootlegged, de formellt planerade produkter,om de byggs alls, är hundar! "
		-- David E. Lundstrom, "A Few Good Men From Univac", MIT Press, 1987

%
"Att ta ett stort steg framåt, måste du göra en serie ändligförbättringar. "
		-- Donald J. Atwood, General Motors

%
"Vi kommer att begrava dig."
		-- Nikita Kruschev

%
"Nu här är något du verkligen kommer att gilla!"
		-- Rocket J. Squirrel

%
"Hur man gör en miljon dollar: Först får en miljon dollar."
		-- Steve Martin

%
"Språk formar vårt sätt att tänka, och bestämmer vad vi kan tänka på."
		-- B. L. Whorf

%
Språket ger en programmerare med en uppsättning av begreppsliga verktyg; om dessa ärotillräcklig för uppgiften, kommer de helt enkelt ignoreras. Till exempel, på allvarbegränsa begreppet pekare tvingar helt enkelt programmeraren att använda envektor plus heltalsaritmetik att genomföra strukturer, pekare, etc. Brautformning och frånvaron av fel kan inte garanteras enbart genom språkfunktioner.
		-- Bjarne Stroustrup, "The C++ Programming Language"

%
"För kärleken av slem ... en dum vägg döds strålar. Hur klibbig kan ya få?"
		-- Post Brothers comics

%
"Byråkrati är fiende till innovation."
		-- Mark Shepherd, former President and CEO of Texas Instruments

%
"En organisation torkar upp om du inte utmana den med tillväxt."
		-- Mark Shepherd, former President and CEO of Texas Instruments

%
"Jag har sett det. Det är skräp."
		-- Marvin the Paranoid Android

%
Vår verksamhet drivs på förtroende. Vi litar på att du betalar i förskott.
		-- Marvin the Paranoid Android

%
"Otrogna i alla åldrar har kämpat för rätten till människa, och har hela tidenvarit orädda förespråkare för frihet och rättvisa. "
		-- Robert Green Ingersoll

%
Historien om uppkomsten av kristendomen har allt att göra med politik,kultur och mänskliga svagheter och ingenting att göra med övernaturliga manipulationav händelser. Hade gudomligt ingripande varit ledstjärnan, säkert tvåårtusenden efter Jesu födelse han inte skulle ha en värld där detfinns fler muslimer än katoliker, mer hinduer än protestanter, och mernontheists än katoliker och protestanter tillsammans.
		-- John K. Naland, "The First Easter", Free Inquiry magazine, Vol. 8, No. 2

%
Jag tycker att du saknar tro på den fjärde dithturbing.
		-- Darse ("Darth") Vader

%
"Alla biblar är konstgjorda."
		-- Thomas Edison

%
"Spock, såg du ser på deras ansikten?""Ja, kapten, en slags ledig belåtenhet."
		-- Thomas Edison

%
"Triumf frihet anarki är nästan (historiskt sett) påhand ... * om * vi kan hålla vänster från att sälja oss som slavar ochRätt från att blåsa upp oss för, säg, de kommande tjugo åren. "
		-- Eric Rayman, usenet guy, about nanotechnology

%
"Gravitation kan inte hållas ansvarig för människor som faller i kärlek."
		-- Albert Einstein

%
"Jag tror att Michael är som lackmuspapper - han alltid försöker att lära sig."
		-- Elizabeth Taylor, absurd non-sequitir about Michael Jackson

%
Även om det inte kan bevisas i efterhand att någon erfarenhet av bollinnehavet,konvertering, uppenbarelse, eller gudomlig extas var bara ett epileptiskt urladdning,vi måste fråga hur man skiljer "verklig transcendens" från neuropatiersom producerar samma extrema realness, djup, ineffability och känslakosmiska enhet. När konton plötsliga konvertering i TLE[Temporal-loben epileptiker] läggs tillsammans med epiphanous uppenbarelserden religiösa traditionen, är paralleller slående. Samma sak gäller för densenaste tidens påstådda UFO bortförda. Sparsamhet ensam argumenterar mot åberoparandar, demoner, eller utomjordingar när naturliga orsaker räcker.- Barry L. Beyerstein, "neuropatologi och Legacy of Spiritual   Besittning ", The Skeptical Inquirer, Vol. XII, nr 3, sid. 255
		-- Elizabeth Taylor, absurd non-sequitir about Michael Jackson

%
"Ett muntligt avtal är inte värt papperet det är tryckt på."
		-- Samuel Goldwyn

%
"Vi ska nå allt större plattityder av prestation."
		-- Richard J. Daley

%
"Med melass du fånga flugor, med vinäger du fånga ingen."
		-- Baltimore City Councilman Dominic DiPietro

%
"Led oss ​​i några ord tyst bön."
		-- Bill Peterson, former Houston Oiler football coach

%
"Jag kunde inte komma ihåg saker tills jag tog att Sam Carnegie kurs."
		-- Bill Peterson, former Houston Oiler football coach

%
"Just nu känner jag att jag har mina fötter på marken så långt som mitt huvudär bekymrad."
		-- Baseball pitcher Bo Belinsky

%
"Nittio procent av baseball är halv mental."
		-- Yogi Berra

%
Två saker är säkra om vetenskap. Det står inte stilla för länge,och det är aldrig tråkigt. Åh, bland några stackars själar, inklusive ävenintellektuella i områden med hög stipendium, är vetenskapen oftamissförståtts. Många ser det som bara en kropp av fakta, som utfärdades frånpå hög måste, obegripliga läroböcker, en samling av oföränderligföreskrifter varas med auktoritära kraft. Andra ser det som ingentingmen en kall, torr smal, grubblande, regelbundet process - den vetenskapligametod: INSKRÄNKT, linjär och vänster brained.Dessa människor är offer för sina egna stereotyper. Dom äravsedd att visa den vetenskapliga världen med en uppsättning skygglappar. Devet ingenting om tumultet, kakofonin, rambunctiousness, ochtendentiousness av den faktiska vetenskapliga processen, än mindrekreativitet, passion och upptäckarglädje. Och det är troligt attvet lite av den ständiga procession av nya insikter och upptäckteratt varje dag, på något sätt, ändra vår uppfattning (om inte deras) avNaturlig värld.- Kendrick Frazier "The Year i Science: En översikt" i   1988 årsbok för vetenskap och framtiden, Encyclopaedia Britannica, Inc.
		-- Yogi Berra

%
"Jackpot: du kan ha en onödig förändring record"
		-- message from "diff"

%
"En advokat kan stjäla mer än hundra män med vapen."
		-- The Godfather

%
Vad är skillnaden mellan en dator försäljare och en bilförsäljare?En bilförsäljare vet när han ljuger.
		-- The Godfather

%
"De som kommer att kunna erövra programvara kommer att kunna erövravärld."
		-- Tadahiro Sekimoto, president, NEC Corp.

%
"Det finns några bra människor i det, men orkestern som helhet är motsvarandetill ett gäng böjd på förstörelse. "
		-- John Cage, composer

%
"Jag tror att användningen av buller att göra musik kommer att öka tills vi når enmusik produceras genom hjälp av elektriska instrument som kommer att göraför musikaliska ändamål som helst och alla ljud som kan höras. "
		-- composer John Cage, 1937

%
Jag gjorde avbryta en prestanda i Holland där de trodde att min musik var så lättatt de inte repetera alls. Och så den första gången när jag fann att ut,Jag repeterade orkestern själv framför publik på 3000 personer ochnästa dag jag repeterade genom den andra satsen - var detta stycke_ Billiga Imitation_ - och de sedan skämdes. Det nederländska folket skämdesoch de uppmanade mig att komma till Holland festivalen och de lovade attrepetera. Och när jag kom till Amsterdam de hade ändrats orkestern, ochigen, hade de inte repeterat. Så de var inte mer förberedd för andra gångenän de hade varit det första. Jag gav dem en föreläsning och berättade för dem att avbrytauppträdandet; De sade sedan över radion att jag hade insisterat på derasavbryta prestanda eftersom de var "otillräckligt Zen."Kan du tro det?
		-- composer John Cage, "Electronic Musician" magazine, March 88, pg. 89

%
"En dag vaknade jag och upptäckte att jag var kär i magar."
		-- Tom Anderson

%
"De flesta människor vill bli befriade från frestelse men skulle vilja att hålla kontakten. "
		-- Robert Orben

%
Regeln om att överleva som en programchef är att ge dem ett nummer ellerge dem ett datum, men aldrig ge dem båda på en gång.
		-- Robert Orben

%
En optimist tror vi lever i den bästa världen möjliga;pessimist fruktar detta är sant.
		-- Robert Orben

%
"Om John Madden steg utanför den 2 februari, tittar ner, och inte se hansfötter, kommer vi att ha ytterligare 6 veckor Pro fotboll. "
		-- Chuck Newcombe

%
Död? Ingen ursäkt för att lägga ut arbete.
		-- Chuck Newcombe

%
Led mig inte in i frestelse ... jag kan hitta det själv.
		-- Chuck Newcombe

%
"När folk är minst säker, de är ofta mest dogmatiska."
		-- John Kenneth Galbraith

%
"Naturen är mycket oamerikansk. Natur aldrig skyndar."
		-- William George Jordan

%
"Vi lär oss av historien som vi lär ingenting av historien."
		-- George Bernard Shaw

%
"Smicker är okej - om du inte andas."
		-- Adlai Stevenson

%
"Konsekvens kräver att du vara så okunnig i dag som du var för ett år sedan."
		-- Bernard Berenson

%
"Toppmöten tenderar att vara som panda parningar. Förväntningarna är alltidhög, och resultaten oftast en besvikelse. "
		-- Robert Orben

%
"Ett stort antal människor tror att de tänker när de bara ordnaderas fördomar. "
		-- William James

%
"Berätta sanningen och springa."
		-- Yugoslav proverb

%
"Den bästa index till en persons karaktär är a) hur han behandlar människor som inte kangör honom något gott och b) hur han behandlar människor som inte kan slå tillbaka. "
		-- Abigail Van Buren

%
"Never inse fakta, om du gör det kommer du aldrig få upp på morgonen."
		-- Marlo Thomas

%
"Livet är ett plagg som vi ständigt ändra, men som aldrig verkar passa."
		-- David McCord

%
"Värdet av äktenskap är inte att vuxna producera barn, men att barnproducera vuxna. "
		-- Peter De Vries

%
"Det är lättare att slåss för principer än att leva upp till dem."
		-- Alfred Adler

%
"Säkerhet är oftast en vidskepelse. Det existerar inte i naturen ... Livet ärantingen ett vågat äventyr eller ingenting. "
		-- Helen Keller

%
"Den som förbinder sig att ställa sig upp som en domare av sanning och kunskap ärskeppsbrutna av skratt av gudarna. "
		-- Albert Einstein

%
"Framgång omfattar en mängd misstag."
		-- George Bernard Shaw

%
"Märket av en omogen man är att han vill dö ädelt för en sak, medanmärket för en mogen man är att han vill leva ödmjukt för en. "
		-- William Stekel

%
"Ja, och jag tycker illa om rendering deras onyttiga carci i dogfood ..."
		-- Badger comics

%
"Är det verkligen du, Fuzz, eller är det Memorex, eller är det strålsjuka?"
		-- Sonic Disruptors comics

%
"De flesta av oss, när allt är sagt och gjort, liksom vad vi vill och späd skälför det efteråt. "
		-- Soren F. Petersen

%
"Du är en varelse av natten, Michael. Wait'll Mamma hör om detta."
		-- from the movie "The Lost Boys"

%
"Plastic pistol. Genialt. Mer kaffe, tack."
		-- The Phantom comics

%
Spelet livet är ett spel av bumeranger. Våra tankar, handlingar och ordtillbaka till oss förr eller senare med häpnadsväckande precision.
		-- The Phantom comics

%
Om först du inte lyckas, kör du om genomsnittet.
		-- The Phantom comics

%
"Ett barn är en person som inte kan förstå varför någon skulle ge bort enhelt bra kattunge. "
		-- Doug Larson

%
"Problemet med att göra något rätt första gången är att ingenuppskattar hur svårt det var. "
		-- Walt West

%
"Tyst tacksamhet är inte mycket nytta för någon."
		-- G. B. Stearn

%
"I principfrågor, stå som en sten, i fråga om smak, simma mednuvarande."
		-- Thomas Jefferson

%
Det första tecknet på mognad är upptäckten att volymratten vänder ocksåvänster.
		-- Thomas Jefferson

%
"Men detta går till elva."
		-- Nigel Tufnel

%
"Gått igenom helvetet? Whaddya föra tillbaka för mig?"
		-- A. Brilliant

%
"Jag vet inte vad deras gripe är. En kritiker är helt enkelt någon som betalas till återge åsikter lättvindigt. ""Kritiker är grinks ochgroinks. "
		-- Baron and Badger, from Badger comics

%
"Jag har fått några amyls. Vi kunde endera parten senare eller, som börjar sitt hjärta."
		-- "Cheech and Chong's Next Movie"

%
"Israel meddelade idag att man ger upp. Den sionistiska staten löseri två veckor, och dess medborgare kommer att sprida till olika utväg samhällenrunt världen. Sade statsminister Yitzhak Shamir, "Vem behöverförvärrande?'"
		-- Dennis Miller, "Saturday Night Live" News

%
"Och, naturligtvis, har du reklamfilmerna där kunniga företagare få ett försprånggenom att använda sina Macintosh-datorer för att skapa den ultimata amerikansk affärsprodukt: en riktigt skarp utseende rapport ".
		-- Dave Barry

%
Handla eller DÖ, människor på jorden![Erbjudande tomrum där det är förbjudet]
		-- Capitalists from outer space, from Justice League Int'l comics

%
"Roman Polanski gör sitt eget blod Han är smart -.. Det är därför hans filmer fungerar"
		-- A brilliant director at "Frank's Place"

%
"Följande är inte för de svaga i hjärtat eller fundamentalister."
		-- Dave Barry

%
"Jag tar honom handla med mig. Jag säger," OK, Jesus, hjälp mig att hitta en bra affär ""
		-- Tammy Faye Bakker

%
Gary Hart: levande bevis på att du * kan * skruva din hjärna ut.
		-- Tammy Faye Bakker

%
Välsignad vara de som initiera livliga diskussioner med hopplöst stum,de skall känna som tandläkare.
		-- Tammy Faye Bakker

%
"Jag tror inte på svepande social förändring manifesteras av en person,om han har en atom vapen. "
		-- Howard Chaykin

%
"Ända fritt klättrade tusen fot vertikal klippa med 60 pounds av redskapfastspänd på din rumpa? "   "Nej.""" Självklart har du inte, du frukt-loop lilla nörd. "- The Mountain Man, en av Dana Carvey: s SNL tecken[dito]
		-- Howard Chaykin

%
"Jag menar, som jag just läst din artikel i lag recept Yale, på sök ochbeslag. Man, var det verkligen där ute. "   "Jag var så HAVERERAD när jag skrev det ..."
		-- John Lovitz, as ex-Supreme Court nominee Alan Ginsburg, on SNL

%
"Hej, jag är professor Alan Ginsburg ... Men du kan kalla mig ... kapten Toke."
		-- John Lovitz, as ex-Supreme Court nominee Alan Ginsburg, on SNL

%
Det är bra att vara smart "för då du vet saker.
		-- John Lovitz, as ex-Supreme Court nominee Alan Ginsburg, on SNL

%
"Tid är pengar och pengar kan inte köpa du älskar och jag älskar din outfit"
		-- T.H.U.N.D.E.R. #1

%
"Kan du inte bara gest hypnotiskt och få honom att försvinna?"    "Det fungerar inte på det sättet. KÖR!"
		-- Hadji on metaphyics and Mandrake in "Johnny Quest"

%
"Du ska inte göra min brödrost arg."
		-- Household security explained in "Johnny Quest"

%
 "Någon har varit elak mot dig! Säg mig vem det är, så jag kan slå honom smakfullt."
		-- Ralph Bakshi's Mighty Mouse

%
"Och barnen ... lära sig något från Susie och Eddie. Om du tror att det finns en maniskt psyko nörd i källare:    1) inte ge honom en chans att träffa dig påhuvudet med en yxa!    2) Fly lokaler ... även om du är i dinunderkläder.    3) varna grannarna och ringa polisen. Men vad du gör ... INTE gå ner på DAMN källaren! "
		-- Saturday Night Live meets Friday the 13th

%
Seger eller nederlag!
		-- Saturday Night Live meets Friday the 13th

%
"Envar har rätt till en * informerade * åsikt."
		-- Harlan Ellison

%
"Det är gardiner för dig,! Pistolen är Mighty Mouse så futuristiska att även* I * vet inte hur det fungerar! "
		-- from Ralph Bakshi's Mighty Mouse

%
"Må de onda krafterna blir förvirrad på vägen till ditt hus."
		-- George Carlin

%
En universitetsfakultet är 500 egoister med gemensam parkering problem.
		-- George Carlin

%
   "Pappa, pappa, gör    Santa Claus försvinna! ""Jag kan inte, son;han blivit förkraftfull. "				     "HO HO HO!"
		-- Duck's Breath Mystery Theatre

%
"Om det inte är högt, fungerar det inte!"
		-- Blank Reg, from "Max Headroom"

%
"Kom ihåg barn, om det finns ett laddat vapen i rummet, vara säker på att du ären hålla den "
		-- Captain Combat

%
Delta: Vi gör aldrig samma misstag tre gånger. - David Letterman
		-- Captain Combat

%
Delta: En riktig man landar där han vill. - David Letterman
		-- Captain Combat

%
Delta: Barnen kommer att älska våra uppblåsbara rutschbanor. - David Letterman
		-- Captain Combat

%
Delta: Vi är Amtrak med vingar. - David Letterman
		-- Captain Combat

%
"Där humor är oroad finns det inga normer - ingen kan säga vad som ärbra eller dåligt, men du kan vara säker på att alla kommer.
		-- John Kenneth Galbraith

%
"Hej igen, Peabody här ..."
		-- Mister Peabody

%
"Det är det bästa sedan professionella golfare på" Ludes. "
		-- Rick Obidiah

%
"Till vänster är marinan där flera höga skåp tjänstemän hålla lyxyachter för weekendkryssningar på Potomac. Några av dessa fartyg är upp till 100fot i längd; Presidentens yacht är över 200 fot i längd, och kanförblir nedsänkt i upp till tre veckor. "
		-- Garrison Keillor

%
"Nå, är social relevans en schtick, som mysterier, social relevans,science fiction..."
		-- Art Spiegelman

%
"Ett av de problem jag har alltid haft med propaganda broschyrer är att de ärverklig tråkigt att titta på. De är bara dåligt utformade. Människor från vänsterofta är mycket välmenande, men de har aldrig haft tid att ta grundkonstruktionklasser, du vet? "
		-- Art Spiegelman

%
"Om du tog alla som någonsin varit i en död visar och ställde upp dem, de skulle sträcka halvvägs till månen och tillbaka ... och ingen av dem skulle vara klaga. "
		-- a local Deadhead in the Seattle Times

%
"Och kom ihåg: onda kommer alltid att segra, eftersom Bra är dum."
		-- Spaceballs

%
Varför är många forskare som använder advokater för medicinskexperiment i stället för råttor?a) Det finns fler advokater än råttor.b) vetenskapsmannens inte blir så emotionellt fäst vid dem.c) Det finns några saker att även råttorkommer inte att göra för pengarna.
		-- Spaceballs

%
"Under loppetVi kan äta din damm,Men när du uppgraderar,Du kommer att arbeta för oss. "
		-- Reed College cheer

%
Pohl lag:Ingenting är så bra att någon, någonstans, kommer inte hata det.
		-- Reed College cheer

%
Pig: Ett djur (Porcus allätare) nära allierad med den mänskliga rasen avprakt och livlighet av dess aptit, vilket emellertid är underlägsen i omfattning,för det balkar på gris.
		-- Ambrose Bierce

%
"Vi har inte för att skydda miljön -. Andra ankomst är nära"
		-- James Watt

%
"Jag tror att Ronald Reagan dag kommer att göra detta land vad det en gång var ... en arktiska vildmarken. "
		-- Steve Martin

%
"Till dig jag en ateist, till Gud, jag är lojal opposition."
		-- Woody Allen

%
Noncombatant: En död Quaker.
		-- Ambrose Bierce

%
"Det finns bara ett sätt att få ett lyckligt äktenskap och så fort jag lära sig vad detär jag gifta igen. "
		-- Clint Eastwood

%
Många människor jag känner tror på positivt tänkande, och så gör I.Jag tror att allt positivt stinker.
		-- Lew Col

%
F: Hur många IBM CPU tar det att utföra ett jobb?A: Fyra; tre för att hålla ner det, och en att slita sitt huvud.
		-- Lew Col

%
Diplomati är konsten att säga "nice doggy" tills du hittar en sten.
		-- Lew Col

%
Harrisberger fjärde lag Lab:Upplevelse är direkt proportionell motmängden utrustning som förstörd.
		-- Lew Col

%
Kapten Penny lag:Du kan lura alla människor en del av dentid, och några av dem alla itid, men du kan inte lura mamma.
		-- Lew Col

%
"För att han är en karaktär som är ute efter sin egen identitet, [He-Man är]en intressant roll för en skådespelare. "
		-- Dolph Lundgren, "actor"

%
"Om Jesus kom tillbaka idag, och såg vad som pågick i hans namn, skulle han aldrigsluta kasta upp. "
		-- Max Von Sydow's character in "Hannah and Her Sisters"

%
"Nietzsche säger att vi kommer att leva samma liv, om och om igen.Gud - Jag måste sitta igenom isen Capades igen ".
		-- Woody Allen's character in "Hannah and Her Sisters"

%
"När det gäller Oral Roberts påstående att Gud sa till honom att han skulle dö om han inte fick $ 20.000.000 av mars, har Guds advokater uppgav att deras klient har inte talat med Roberts under flera år. Off the record, har Gud förklarat att "Om jag hade velat is lilla padda, skulle jag ha gjort det för länge sedan."
		-- Dennis Miller, SNL News

%
"Endast hycklare är verkligen ruttet till kärnan."
		-- Hannah Arendt.

%
Quod licet Iovi non licet Bovi.(Vad Jove kan göra, inte är tillåtet att en ko.)
		-- Hannah Arendt.

%
"Jag misstror en man som säger" när ". Om han måste vara noga med att inte dricka förmycket, beror det på att han inte är att lita på när han gör. "
		-- Sidney Greenstreet, _The Maltese Falcon_

%
"Jag misstror en nära mun man. Han plockar generellt fel tid att prataoch säger fel saker. Talking är något du inte kan göra klokt,om du håller i praktiken. Nu, sir, kommer vi att tala om du vill. Jag ska berättadu rätt ut, jag är en man som gillar att prata med en man som gillar att prata. "
		-- Sidney Greenstreet, _The Maltese Falcon_

%
Alla extremister ska tas ut och sköt.
		-- Sidney Greenstreet, _The Maltese Falcon_

%
"Sextiotalet var bra för dig, inte de?"
		-- George Carlin

%
"Stanna här, Audrey - detta är mellan mig och grönsaker!"
		-- Seymour, from _Little Shop Of Horrors_

%
Från skarpa hjärnor kommit ... pekade huvuden.
		-- Bryan Sparrowhawk

%
Det finns två typer av egoister: 1) De som medger det 2) Resten av oss
		-- Bryan Sparrowhawk

%
"Bilden är ganska dystra, herrar ... Världens klimat förändras,däggdjuren tar över, och vi alla har en hjärna ungefär lika stor som envalnöt."
		-- some dinosaurs from The Far Side, by Gary Larson

%
"Vi amerikaner, vi är en enkel folk ... men pissa oss, och vi kommer att bombadina städer. "
		-- Robin Williams, _Good Morning Vietnam_

%
Varför inte hajar äta advokater? Professionell artighet.
		-- Robin Williams, _Good Morning Vietnam_

%
"Du vet, vi har vunnit priser för denna skit."
		-- David Letterman

%
Det var synd stannade handen."Synd att jag inte har några fler kulor," tänkte Frito.
		-- _Bored_of_the_Rings_, a Harvard Lampoon parody of Tolkein

%
En bra USENET motto skulle vara: en. "Tillsammans en stark gemenskap." b. "Datorer R Us." c. "Jag är trött på programmering, jag tror jag ska bara skruva runt ett tag på     företagets tid. "
		-- A Sane Man

%
"Han inte köra för omval. 'Politik tar dig i kontakt med allapersoner som du skulle ge vad som helst för att undvika, sade han. 'Jag stannar hemma. "
		-- Garrison Keillor, _Lake_Wobegone_Days_

%
"Om du levt i dag som om det vore din sista, skulle du köpa upp en låda med raketer ochavfyra dem alla, skulle inte du? "
		-- Garrison Keillor

%
"Mr Spock dukar till en kraftfull parning lust och nästan dödar kapten Kirk."
		-- TV Guide, describing the Star Trek episode _Amok_Time_

%
"Dålig människa ... han var som en anställd till mig."
		-- The police commissioner on "Sledge Hammer" laments the death of his bodyguard

%
"Tro mig. Jag vet vad jag gör."
		-- Sledge Hammer

%
"Hej. Det här är Dan Cassidy telefonsvarare. Lämna ditt namn ochantal ... och efter att jag har manipulerat bandet, kommer ditt meddelande implicerade dig i ett federalt brott och att uppmärksammas av F.B.I ... BEEEP "
		-- Blue Devil comics

%
"Alla Guds barn är inte vacker. De flesta av Guds barn är i själva verket,knappt presentabel. "
		-- Fran Lebowitz

%
"Om sanningen är skönhet, hur kommer ingen har sitt hår gjort i biblioteket?"
		-- Lily Tomlin

%
Som gudarna skulle förstöra de först lära BASIC.
		-- Lily Tomlin

%
"Titta! Där! Evil! .. Ren och enkel, total ondska från åttonde dimensionen!"
		-- Buckaroo Banzai

%
"Jag kan vara syntetiska, men jag är inte dum"
		-- the artificial person, from _Aliens_

%
"Det enda sättet jag kan förlora detta val är om jag fångad i sängen med en dödflicka eller en levande pojke. "
		-- Louisiana governor Edwin Edwards

%
David Letterman s "Saker som vi kan vara stolta över som amerikaner":* Största antalet medborgare som faktiskt har bordade ett UFO* Många tidningar funktionen "RÖRA"* timma motell* De allra flesta Elvis filmer görs här* Inte bara ge upp direkt under andra världskriget som en delländer som vi skulle kunna nämna* Goatees & Van Dykes tros endast bäras av weenies* Våra skötsam golfproffs* Fabulous babes kust till kust
		-- Louisiana governor Edwin Edwards

%
"Fara, har du inte sett det sista av mig!"   "Nej, men det första ni vänder min mage!"
		-- The Firesign Theatre's Nick Danger

%
Ber till Gud, men hålla rodd till stranden.
		-- Russian Proverb

%
"Oroa dig inte om folk stjäl dina idéer. Om dina idéer är något bra,du måste ramma dem ner folks halsar. "
		-- Howard Aiken

%
"När någon säger 'teoretiskt," de egentligen menar `inte riktigt."
		-- David Parnas

%
"Inga problem är så formidabel att du inte kan gå ifrån det."
		-- C. Schulz

%
"Den goda kristna ska akta sig för matematiker och alla dem som görtomma profetior. Faran finns redan att matematiker har gjortett förbund med djävulen mörkare anda och begränsa man iobligationer i helvetet. "
		-- Saint Augustine

%
"För mannen som har allt ... Penicillin."
		-- F. Borquin

%
 "Jag har äntligen lärt sig vad` uppåt kompatibla "betyder. Det betyder att vi  får behålla alla våra gamla misstag. "
		-- Dennie van Tassel

%
"Sättet att världen är att prisa döda helgon och åtala levande sådana."
		-- Nathaniel Howe

%
"Det är en hund-äta-hundvärlden där ute, och jag bär Milkbone ware."
		-- Norm, from _Cheers_

%
En gång på en tillställning, sade Gladstone till Disraeli, "Jag förutspår, Sir, attdu kommer att dö antingen genom hängning eller någon vile sjukdom ". Disraeli svarade"Det beror, Sir, på om jag omfamna era principer eller dinhusmor."
		-- Norm, from _Cheers_

%
"Han vet inte mig vewy väl, DO han?" - Bugs Bunny
		-- Norm, from _Cheers_

%
"Jag ska råna att rik person och ge den till någon fattig förtjänar slusk. Det kommer * bevisa * Jag är Robin Hood. "
		-- Daffy Duck, Looney Tunes, _Robin Hood Daffy_

%
"Skulle jag slå på gasen om min kompis Mugsy var där?"   "Du kanske, kanin, kanske du!"
		-- Looney Tunes, Bugs and Thugs (1954, Friz Freleng)

%
"Consequences, Schmonsequences, så länge jag är rik."
		-- Looney Tunes, Ali Baba Bunny (1957, Chuck Jones)

%
"Och tror du (FOP att jag) att jag kunde vara Scarlet pumpernickel?"
		-- Looney Tunes, The Scarlet Pumpernickel (1950, Chuck Jones)

%
"Nu har jag pärlan på dig med min sönderfallande pistol. Och när detupplöses, sönderdelas det. (Drar utlöser) Nå, vad du vet,det upplöstes. "
		-- Duck Dodgers in the 24th and a half century

%
"Döda Wabbit, döda Wabbit, Döda Wabbit!"
		-- Looney Tunes, "What's Opera Doc?" (1957, Chuck Jones)

%
"Jag vill dina pengar, eftersom Gud vill ha dina pengar!"
		-- The Reverend Jimmy, from _Repo_Man_

%
"Majoriteten av de dumma är oövervinnelig och garanteras för all framtid. Denterror deras tyranni, dock lindras genom deras brist på konsekvens. "
		-- Albert Einstein

%
"Du visa mig en amerikan som kan hålla hans mun och jag ska äta honom."
		-- Newspaperman from Frank Capra's _Meet_John_Doe_

%
"Och vi hörde honom utropaNär han började ströva:'Jag är ett hologram, barn,försök inte detta hemma! "- Bob våld
		-- Howie Chaykin's little animated 3-dimensional darling, Bob Violence

%
"Sovjetunionen, som har klagat nyligen om påstådda antisovjetiskteman i amerikansk reklam, lämnat in en officiell protest denna vecka motFord Motor Companys nya kampanj: 'Hej du stinkande fett ryska, får av min Ford Escort. "
		-- Dennis Miller, Saturday Night Live

%
"Det finns gott hopp om symbolik i det faktum att flaggor inte vågen i ett vakuum."
		-- Arthur C. Clarke

%
"De borde göra stum smaksatt kattmat." --Gallagher
		-- Arthur C. Clarke

%
"Inte bara är Gud död, men bara försöka hitta en rörmokare på helgerna."
		-- Woody Allen

%
"Klockan är tio ... Vet du var dina AI program?" - Peter Oakley
		-- Woody Allen

%
"Ah, du vet vilken typ. De gillar att skylla allt på judar eller svarta,För om de inte kunde, skulle de behöva vakna upp till det faktum att livet är en stor,skrämmande, strålande, komplex och slutligen outgrundliga crapshoot - och det endaAnledningen till att de inte kan hålla jämna steg är att de är ett gäng misfits och förlorare. "
		-- an analysis of neo-Nazis and such, Badger comics

%
"Intressant undersökning i nuvarande Journal of Abnormal Psychology: New YorkStaden har en högre andel personer som du bör inte göra några plötsliga rörelserrunt än någon annan stad i världen. "
		-- David Letterman

%
"Turister - ha lite kul med New Yorks hårdkokta cabbies När du får.till din destination, säg till din förare, "Betala? jag lifta."
		-- David Letterman

%
"En antropolog vid Tulane har precis kommit tillbaka från en studieresa till NewGuinea med rapporter om en stam så primitivt att de har Tide men intenya Tide med citron-fresh Borax. "
		-- David Letterman

%
"Baserat på vad du vet om honom i historieböckerna, vad tror du AbrahamLincoln skulle göra om han levde idag?1) Att skriva sina memoarer av inbördeskriget.2) Att ge råd ordföranden.3) Desperat clawing vid insidan av hanskista. "
		-- David Letterman

%
"Om Rick Schroder och Gary Coleman hade en kamp på TV med poolköer, vem skulle vinna?1) Rick Schroder2) Gary Coleman3) TV-tittande allmänheten "
		-- David Letterman

%
"Om du börjar tvivla vad jag säger, du är förmodligen hallucinerar. "
		-- The Firesign Theatre, _Everything you know is Wrong_

%
Vad att göra i händelse av en främmande attack:    1) Hide under sätet för din plan och titta bort.    2) Undvik kontakt med ögonen.    3) Om det inte finns några ögon, undvika all kontakt.
		-- The Firesign Theatre, _Everything you know is Wrong_

%
"Kärnvapenkrig skulle verkligen tillbaka kabeln."
		-- Ted Turner

%
"Du tweachewous miscweant!"
		-- Elmer Fudd

%
"Jag såg _Lassie_. Det tog mig fyra visar att räkna ut varför den håriga ungen aldrigeker. Jag menar, han kunde rulla över och allt det där, men det förtjänar en serie? "
		-- the alien guy, in _Explorers_

%
"Öppen kanal D ..."
		-- Napoleon Solo, The Man From U.N.C.L.E.

%
Rädda valarna. Samla hela uppsättningen.
		-- Napoleon Solo, The Man From U.N.C.L.E.

%
Stödja Mental Health. Eller jag ska döda dig.
		-- Napoleon Solo, The Man From U.N.C.L.E.

%
"Pyramiden öppnar!"   "Vilken?""Den med allt större hål i det!"
		-- The Firesign Theatre

%
"Calling J-Man Kink. Ringa J-Man Kink. Hash missil seende, målLos Angeles. Bortse från personliga känslor om staden och avlyssna. "
		-- The Firesign Theatre movie, _J-Men Forever_

%
"Min känsla av mening är borta! Jag har ingen aning om vem jag är!"    "Herregud ... Du har .. Du har gjort honom till en demokrat!"
		-- Doonesbury

%
"Du har fel, du ol 'mässing knäppt fascistiska poop!"
		-- Bloom County

%
"Din mor var en hamster och din far luktade fläderbär!"
		-- Monty Python and the Holy Grail

%
"Väljarna har talat, de jävlarna ..."
		-- unknown

%
"Jag föredrar att tro att Gud är inte död, bara full"
		-- John Huston

%
"Var det. Aloha."
		-- Steve McGarret, _Hawaii Five-Oh_

%
"När det blir konstigt, konstiga tur pro ..."
		-- Hunter S. Thompson

%
"Säg yur böner, yuh lopp Pickin varmint!"
		-- Yosemite Sam

%
"Det ... Jag har kört ringarnas runt du logiskt"
		-- Monty Python's Flying Circus

%
... Veloz är omöjlig att skilja från hundratals andra elektronikföretagi dalen, som drivs av ivriga unga ingenjörer lutad över minnesdumpar sentframåt natten. Skillnaden är att ett gäng själv erkände "bil nötter"tjänar pengar gör vad de älskar: att skriva kod och köra fort.
		-- "Electronics puts its foot on the gas", IEEE Spectrum, May 88

%
"Bara fakta, frun"
		-- Joe Friday

%
"Jag har fem dollar för var och en av er."
		-- Bernhard Goetz

%
Mausoleum: Den sista och roligaste dårskap för de rika.
		-- Ambrose Bierce

%
Rikedom: En gåva från himlen betyda, "Detta är min älskade son, i vilken jagär mycket nöjd. "
		-- John D. Rockefeller, (slander by Ambrose Bierce)

%
Allt är antingen heligt eller profan.Den förstnämnda till ecclesiasts få vinst;Den senare till djävulen appertain.
		-- Dumbo Omohundro

%
Saint: En död syndare reviderad och redigeras.
		-- Ambrose Bierce

%
Fyrtiotvå.
		-- Ambrose Bierce

%
Saktmod: Mindre vanliga tålamod planerar en hämnd som är värt mödan.
		-- Ambrose Bierce

%
Absolut: Oberoende, oansvarigt. En absolut monarki är en i vilkensuveräna gör som han vill så länge han vill mördarna. Intemånga absoluta monarkier är kvar, de flesta av dem har ersatts avbegränsade monarkier, där suveräna makt för ont (och goda) ärkraftigt begränsas, och av republikerna, som styrs av en slump.
		-- Ambrose Bierce

%
Absolutist: En svag person som ger efter för frestelsen att förneka sig själv ennöje. En absolutist är en som avstår från allt, mennedlagd röst, och i synnerhet från inaktivitet i andras angelägenheter.
		-- Ambrose Bierce

%
Alliance: I den internationella politiken, en förening av två tjuvar som har sinhänder så djupt in i varandras ficka som de kan inte separatplundring tredjedel.
		-- Ambrose Bierce

%
Olydnad: Den guldkant till molnet av slaveri.
		-- Ambrose Bierce

%
Egoist: En person med låg smak, mer intresserad av sig själv än i mig.
		-- Ambrose Bierce

%
Administration: En genial abstraktion i politik, som syftar till att ta emotsparkar och manschetter på grund av premier eller president.
		-- Ambrose Bierce

%
En sparad krona är en krona för att slösa.
		-- Ambrose Bierce

%
Ocean: En vattenförekomst som upptar cirka två tredjedelar av en värld för människan -som inte har några gälar.
		-- Ambrose Bierce

%
Läkare: En på vilken vi sätter vårt hopp när sjuk och våra hundar när väl.
		-- Ambrose Bierce

%
Filosofi: En rutt av många vägar som leder från ingenstans till ingenting.
		-- Ambrose Bierce

%
Politik: En strid intressen maskerats som en tävling av principer.Genomförandet av offentliga angelägenheter för privat fördel.
		-- Ambrose Bierce

%
Politiker: En ål i den grundläggande leran på vilken överbyggnadorganiserade samhället föds. När han slingrar han misstag agitationen avsvansen för darrande av byggnaden. Jämfört med statsman,han lider av nackdelen av att vara vid liv.
		-- Ambrose Bierce

%
Be: Att be att universums lagar ogiltigförklaras till förmån för en endaStällaren UPPENBARLIGEN ovärdigt.
		-- Ambrose Bierce

%
Ordförandeskapet: Den smord gris inom omgång amerikansk politik.
		-- Ambrose Bierce

%
Snabel: Den rudimentära organ av en elefant som tjänar honom på platsav kniv och gaffel som Evolution ännu har förnekat honom. för ändamålhumor det populärt kallas en trunk.
		-- Ambrose Bierce

%
"Dagens robotar är mycket primitiva, kapabla att förstå endast ett fåtal enkla instruktioner som "gå till vänster", "gå till höger" och "bygga bil". "
		-- John Sladek

%
"I kampen mellan dig och världen, tillbaka i världen."
		-- Frank Zappa

%
Här är en Appalachian version av ledningens svar till dem som ärberörs av ödet av projektet:"Oroa dig inte mule. Bara ladda vagnen."
		-- Mike Dennison's hillbilly uncle

%
Illa vald abstraktion är särskilt tydligt i utformningen av ADAruntime-system. Gränssnittet till ADA runtime systemet är så opak attdet är omöjligt att modellera eller förutsäga dess prestanda, vilket gör det effektivtvärdelös för realtidssystem. - Marc D. Donner och David H. Jameson.
		-- Mike Dennison's hillbilly uncle

%
"Att mot tortyr borde vara en slags tvåparti sak."
		-- Karl Lehenbauer

%
"Här kommer Bill hund."
		-- Narrator, Saturday Night Live

%
Sex är som luft. Det är bara en stor sak om du inte kan få någon.
		-- Narrator, Saturday Night Live

%
"Ha en medvetenhet om bidrag - till ditt schema, ditt projekt,vårt bolag."
		-- A Group of Employees

%
"Fråga inte vad en grupp anställda kan göra för dig. Men fråga vad kanAlla anställda gör för en grupp anställda. "
		-- Mike Dennison

%
En kväll Mr Rudolph Block, New York, befann sig sittande vid middagentillsammans med Mr Percival Pollard, den framstående kritiker.   "Mr Pollard", sade han, "min bok, _The biografi av en död Cow_, är publicerade anonymt, men du kan knappast vara okunnig om dess författarskap. Ändå att granska det ni talar om det som ett verk av den Idiot av århundradet. Tror du att en rättvis kritik? "   "Jag är mycket ledsen, min herre", svarade kritiker, vänligt ", men det gjorde intefalla mig att du verkligen inte kan önska allmänheten att veta vem som skrev den. "
		-- Ambrose Bierce

%
Många alligatorer kommer att dödas,men träsket förblir.
		-- Ambrose Bierce

%
Vad gudarna skulle förstöra de först underkasta sig en Standards Committee IEEE.
		-- Ambrose Bierce

%
Det är nu. Senare är senare.
		-- Ambrose Bierce

%
"Jag kommer att göra några fynd med hårdvara terrorism."
		-- Peter da Silva

%
"Om jag inte återvänder till talarstolen i helgen, kommer miljontals människor gåråt helvete."
		-- Jimmy Swaggart, 5/20/88

%
"Dump kryddor. Om vi ​​är ätas, behöver vi inte att smaka gott."
		-- "Visionaries" cartoon

%
"Shit, om du gör mig att gråta längre, du dimma upp min hjälm."
		-- "Visionaries" cartoon

%
Jag vill inte vara ung igen, jag vill bara inte att få någon äldre.
		-- "Visionaries" cartoon

%
Vigsel: En otrolig metafysiska bluff för att titta på Gud ochlag som dras in i affärer i din familj.
		-- O. C. Ogilvie

%
  "Nödsituation!" Sgiggs skrek, mata ut sig från badkaret som det varen brinnande bil. "Ring" ett "Få room service! Code Red" Stiggs var påtelefonen omedelbart, beställa mer ros blommar, eftersom det, enligthonom hade de som flyter i badkaret plötsligt förlorat sin lukt. "Jag kräverlukt ", han shrilled." Jag förväntar total oavbruten lukt från dessaf * cking rosor. "  Tyvärr har tjänsten kaptenen inte inse att Stiggs situationeninvolverade femtio rosor. "Vad ska jag göra med det här?" Stiggs sneered påden weaseling hotell goon när han dök upp på vår dörr som innehar en enda blommaflytande i en brandy glas. Stiggs s harang var stor. "Ser du dettabadkar? Märker du någon skillnad mellan storleken på badkaret ochStorleken på den spinkiga bunt kronblad i din hand? Jag behöver total bad täckning.Jag behöver en helt fast skikt av rosor runt mig som bloss fabrikerinne, angriper mig med deras lukt och power-ramma stor stinkandekoncentrationer av ökade lukt mina näsborrar tills jag slösat med glädje. "Det dröjde inte länge innan vi fick så missnöjda med denna inkompetens som vibultad.- Den Helt Monstrous, Mind-Rostning Summer of O.C. och Stiggs,   National Lampoon, oktober 1982
		-- O. C. Ogilvie

%
När den är felaktig, är det, åtminstone * auktoritet * felaktig.
		-- Hitchiker's Guide To The Galaxy

%
Vi beslutade att det var natten igen, så vi slog läger i tjugo minuter och drackytterligare sex öl på en ung Life campingplats. O.C. kom in i tillsynsvuxnes sovsäck och sprang runt i den. "Detta är domens dag och jag ären skrämmande syn ", skrek han. Då värmen O.C. Ralph iväska.- Den Helt Monstrous, Mind-Rostning Summer of O.C. och Stiggs,   National Lampoon, oktober 1982
		-- Hitchiker's Guide To The Galaxy

%
Voodoo Programmering: Saker programmerare gör att de vet inte fungera utande försöker ändå, och som ibland faktiskt fungerar, såsom kompileraallt.
		-- Karl Lehenbauer

%
Detta är naturligtvis att helt oinformerad spekulationer om att jag delta i hjälpastödja mitt fördomar mot sådan inblandning ... men där har du det.- Peter da Silva, spekulera om varför ett datorprogram som hade varitändrats för att göra något som han inte godkänner, inte fungerade
		-- Karl Lehenbauer

%
"Denna kunskap jag fortsätta är den finaste glädje jag någonsin har känt. Jag kundeKnappt ge upp att jag kunde själva luften som jag andas. "
		-- Paolo Uccello, Renaissance artist, discoverer of the laws of perspective

%
"Jag fick alla att betala upp framför ... då jag sprängde deras planet."  "Nu varför inte jag tänker på det?"
		-- Post Bros. Comics

%
"Atomic batterier till makten, turbiner för att påskynda."
		-- Robin, The Boy Wonder

%
F-15 Eagle:Om det är det, vi skjuter det ner. Om det är nere, vi blåsa upp det.
		-- A McDonnell-Douglas ad from a few years ago

%
"Amiga är den enda dator där du kan köra en multitaskingoperativsystem och få realtidsprestanda, out of the box ".
		-- Peter da Silva

%
"Det är min cookie-fil och om jag komma fram till något som är haltande och jag gillar det,det går i. "
		-- karl (Karl Lehenbauer)

%
Att erkänna AT & T Bell Laboratories för företagens innovation, för sinUppfinningen av cellulära mobilkommunikation, IEEE president Russell C. Drewhänvisas till den cellulära telefonen som en "grundläggande nödvändighet." Hur gånger harändrats, sade en observatör: många i rummet påminde tillkomsten avdirekt uppringning.
		-- The Institute, July 1988, pg. 11

%
... Sovjet har förmågan att prova stora projekt. Om det finns ett mål,till exempel när Gorbatjov säger att de kommer att ha atomdrivenhangarfartyg, är fallet stängd - det är det. De kommer att koncentrerapå problemet, gör ett dåligt jobb, och senare betala priset. De verkligen intebry sig om vad priset är.- Viktor Belenko, MiG-25 stridspilot som hoppade av 1976   "Defense Electronics", vol 20, nr 6, sid. 100
		-- The Institute, July 1988, pg. 11

%
Det är något du måste förstå om det sovjetiska systemet. De har denförmåga att koncentrera alla sina ansträngningar på en viss design och utveckla allakomponenter samtidigt, men ibland utan riktig testning. Då de slutarmed en teknisk katastrof som Tu-144. I en teknik lopp påtiden, att flygplanet var två månader före Concorde. Fyra Tu-144Sbyggdes; två har kraschat, och två är i museer. Concorde har varitflygande säkert i över 10 år.- Viktor Belenko, MiG-25 stridspilot som hoppade av 1976   "Defense Electronics", vol 20, nr 6, sid. 100
		-- The Institute, July 1988, pg. 11

%
DE: Sovjet verkar ha svårt att genomföra modern teknik.     Vill du kommentera det?Belenko: Tja, låt oss tala om flygmotor livstid. När jag flögMiG-25, dess motorer hade en total livslängd på 250 timmar.DE: Är det medeltid mellan-fel?Belenko: Nej, motorn är klar; den skrotas.DE: Du menar att de dra ut och kasta bort det, inte ens se över det?Belenko: Det är korrekt. Översyn är för dyrt.DE: Det är absurt låg av fria internationella standarder.Belenko: Jag vet.- En intervju med Viktor Belenko, MiG-25 stridspilot som hoppade av 1976   "Defense Electronics", vol 20, nr 6, sid. 102
		-- The Institute, July 1988, pg. 11

%
"Jag har en vän som precis kommit tillbaka från Sovjetunionen, och berättade människorDet är hungriga för information om väst. Han tillfrågades om mångasaker, men jag kommer att ge dig två exempel som är mycket avslöjande om livet iSovjetunionen. Den första frågan han tillfrågades var om vi hade exploderandeTV-apparater. Du ser, de har ett problem med bildrör på färgTV-apparater, och många exploderar. De trodde vi måste haproblem med dem också. Den andra frågan han tillfrågades ofta var därförCIA hade dödat Samantha Smith, den lilla flickan som besökte Sovjetunionen ennågra år sedan; deras propaganda är mycket effektiv.- Viktor Belenko, MiG-25 stridspilot som hoppade av 1976   "Defense Electronics", vol 20, nr 6, sid. 100
		-- The Institute, July 1988, pg. 11

%
"... Jag skulle kunna godta denna öppenhet, glasnost, perestrojka, eller vad du villatt kalla det om de gjorde dessa saker: avskaffa ett partisystem; öppnaSovjetiska gränsen och låta sovjetiska folket att resa fritt; tillåta den sovjetiskamänniskor att få verklig fri företagsamhet; låta västerländska affärsmän att göra affärerdär, och tillåta yttrandefrihet och pressen. Men än så länge, helaLandet är som ett koncentrationsläger. Taggtråden på staketet runtSovjetunionen är att hålla folk inne i mörkret. Denna öppenhet somdu ser, alla dessa förändringar, är kosmetiska och de har utformatsatt imponera kortsynta, naiva, ibland dumma västerländska ledare. Dessaledare forsa över Gorbatjov, i hopp om att göra affärer med Sovjetunionen ellerblidka den. Han kommer att säga: "Ja, vi kan göra affärer!" Detta medan hansmilitär maskin i Afghanistan har dödat över en miljon människor ur enbefolkning på 17 miljoner. Kan ni föreställa er det?- Viktor Belenko, MiG-25 stridspilot som hoppade av 1976   "Defense Electronics", vol 20, nr 6, sid. 110
		-- The Institute, July 1988, pg. 11

%
"Kom ihåg Kruschev: han försökte göra alltför många saker för fort, och han varavlägsnas i onåd. Om Gorbatjov försöker förstöra systemet eller göra alltförmånga grundläggande förändringar av det, tror jag att systemet kommer att bli av med honom.Jag är inte en statsvetare, men jag förstår systemet mycket väl.Jag tror att han kommer att ha en "hjärtattack" eller går i pension eller tas bort. Han ärupp mot en tegelvägg. Om du tror att de kommer att ändra allt ochbli en fri, öppet samhälle, glöm det! "- Viktor Belenko, MiG-25 stridspilot som hoppade av 1976   "Defense Electronics", vol 20, nr 6, sid. 110
		-- The Institute, July 1988, pg. 11

%
FORTRAN? Den syntaktiskt felaktiga uttalande "DO 10 I = 1,10" kommer att tolka ochgenerera kod skapa en variabel, DO10I, enligt följande: "DO10I = 1,10" Om detinte skrämma dig, bör det.
		-- The Institute, July 1988, pg. 11

%
"Jag visste då (1970) att en 4-kbyte minidator skulle kosta så mycket somett hus. Så jag resonerade att efter college, skulle jag behöva leva billigt ien lägenhet och lägga alla mina pengar till att äga en dator. "
		-- Apple co-founder Steve Wozniak, EE Times, June 6, 1988, pg 45

%
HP hade en unik policy att låta sina ingenjörer att ta delar från lager somlänge de byggde något. "De tänkte att med varje design, var defå en bättre ingenjör. Det är en politik som jag uppmanar alla företag att anta. "- Apples grundare Steve Wozniak, "Will Wozniak klass ger Apple till lärare?"   EE Times den 6 juni 1988, pg 45
		-- Apple co-founder Steve Wozniak, EE Times, June 6, 1988, pg 45

%
"Jag vill bara vara en bra ingenjör."- Steve Wozniak, en av grundarna av Apple Computer, ingå sitt inledningsanförande   vid 1988 AppleFest
		-- Apple co-founder Steve Wozniak, EE Times, June 6, 1988, pg 45

%
"Det har alltid varit Babels torn slags käbbel i Unix, men dettaär den mest extrema formen någonsin. Detta innebär åtminstone flera år av förvirring. "- Bill Gates, grundare och ordförande i Microsoft,   om Open Systems Foundation
		-- Apple co-founder Steve Wozniak, EE Times, June 6, 1988, pg 45

%
"När du är osäker, skriva ut dem."
		-- Karl's Programming Proverb 0x7

%
"Om du vill ha de bästa saker att hända i företagens liv du måste hitta sättatt vara öppen för den ovanliga personen. Du får inte innovation som endemokratiska processen. Du får nästan det som en anti-demokratisk process.Visst får du det som en anthitetical process, så du måste ha enmiljö där kroppen människor är verkligen mottagliga för förändringar och kanhantera de konflikter som uppstår ur förändring en innovation. "- Max DePree, ordförande och VD för Herman Miller Inc.,   "Herman Millers Secrets of Corporate kreativitet",   The Wall Street Journal, 3 maj 1988
		-- Karl's Programming Proverb 0x7

%
"I näringslivet, jag tror att det finns tre viktiga områden vilka avtalkan inte ta itu med, det gäller konflikten området förändringar och området att nåpotential. För mig ett förbund är en relation som bygger på sådana sakersom delade ideal och delade värdesystem och delade idéer och deladeöverenskommelse om de processer som vi kommer att använda för att arbeta tillsammans. Imånga fall utvecklas till verkliga kärleksrelationer. "- Max DePree, ordförande och VD för Herman Miller Inc., "Herman Millers   Secrets of Corporate kreativitet ", The Wall Street Journal, 3 maj 1988
		-- Karl's Programming Proverb 0x7

%
Ett annat mål är att etablera en relation ", där det är OK för allaatt göra sitt bästa. Det finns en väldig massa människor i ledningen som verkligenvill inte underordnade att göra sitt bästa, eftersom det blir att vara myckethotfull. Men vi har funnit att både internt och med utanfördesigners om vi är villiga att ha denna typ av relation och om vi ärvillig att vara utsatta för vad som kommer att komma ut av det, vi får riktigt braarbete."- Max DePree, ordförande och VD för Herman Miller Inc., "Herman Millers   Secrets of Corporate kreativitet ", The Wall Street Journal, 3 maj 1988
		-- Karl's Programming Proverb 0x7

%
I sin bok, berättar Mr DePree historien om hur designern George Nelson uppmanadeatt bolaget tar också på Charles Eames i slutet av 1940-talet. Max far,J. DePree, en av grundarna av bolaget med Herman Miller 1923, frågade MrNelson om han verkligen ville dela de begränsade möjligheterna i en sedan-smallföretag med en annan designer. "George svar var ungefär så här:'Charles Eames är en ovanlig talang. Han är väldigt annorlunda från mig. DeFöretaget behöver oss båda. Jag vill väldigt gärna ha Charles Eames andel ivad potential som finns. ""- Max DePree, ordförande och VD för Herman Miller Inc., "Herman Millers   Secrets of Corporate kreativitet ", The Wall Street Journal, 3 maj 1988
		-- Karl's Programming Proverb 0x7

%
Mr DePree tror deltagande kapitalismen är den våg av framtiden. DeUS arbetskraften, menar han, "fler och fler krav på att ingå ikapitalistiska systemet och om vi inte hitta sätt att få det kapitalistiska systemetatt vara ett inkluderande system snarare än det exklusiva systemet har varit, vi äralla stora problem. Om vi ​​inte hitta sätt att börja förstå attkapitalismens högsta potential ligger i det gemensamma bästa, inte i de enskildabra, då vi riskerar själva systemet. "- Max DePree, ordförande och VD för Herman Miller Inc., "Herman Millers   Secrets of Corporate kreativitet ", The Wall Street Journal, 3 maj 1988
		-- Karl's Programming Proverb 0x7

%
Mr DePree förväntar sig också en "enorm social förändring" på alla arbetsplatser. "NärJag började först arbeta 40 år sedan, var en fabrik handledare fokuserat påprodukt. Idag är det drastiskt annorlunda, på grund av den sociala miljön.Det är inte ovanligt att en arbetstagare att komma fram på sitt skift och har vissa familjenproblem att han inte vet hur man ska lösa. Exemplet jag vilja använda är enkillen som kommer in och säger "detta inte kommer att bli en bra dag för mig, min sonär i fängelse på en berusad körning laddning och jag vet inte hur man skall höja borgen. "Vad det betyder är att om handledaren vill produktivitet, måste han vetahur man skall höja borgen. "- Max DePree, ordförande och VD för Herman Miller Inc., "Herman Millers   Secrets of Corporate kreativitet ", The Wall Street Journal, 3 maj 1988
		-- Karl's Programming Proverb 0x7

%
Dårar ignorera komplexitet. Pragmatiker lida det.Vissa kan undvika det. Genier ta bort den.
		-- Perlis's Programming Proverb #58, SIGPLAN Notices, Sept.  1982

%
"Vad händer om" är ett varumärke som tillhör Hewlett Packard, så sluta använda den i dinmeningar utan tillstånd, eller riskerar att bli stämd.
		-- Perlis's Programming Proverb #58, SIGPLAN Notices, Sept.  1982

%
Nu, om världens ledare - människor som är ledare på grund avpolitiska, militära eller finansiella styrka, och inte nödvändigtvis visdom ellerhänsyn till mänskligheten - om dessa ledare hantera inte att dra ossöver randen till planet självmord, trots att de ibland pompösaförslag som de kan känna sig tvungna att göra det, kan vi överleva bortom1988.
		-- George Rostky, EE Times, June 20, 1988 p. 45

%
De väsentliga idéer Algol 68 var att hela språket bör varapreciseras och att alla bitar ska passa ihop smidigt.Grundtanken bakom Pascal var att det inte spelade någon roll hur vag denspråkspecifikationen var (det tog * år * att klargöra) eller hur många grovakanter fanns, så länge som CDC Pascal kompilatorn var snabb.
		-- Richard A. O'Keefe

%
"Vi kom. Vi såg. Vi sparkade sin röv."
		-- Bill Murray, _Ghostbusters_

%
"Stjärnorna är gjorda av samma atomer som jorden." Jag brukar plocka en litenämne som detta att ge en föreläsning om. Poeter säger vetenskapen tar bort frånskönhet av stjärnorna - bara droppar av gas atomer. Ingenting är "bara". Även jag kanse stjärnorna på en ökennatten, och känner dem. Men ser jag mer eller mindre?Vidden av himlen sträcker min fantasi - fastnat på denna karusellmin lilla ögat kan fånga en miljon år gammal ljus. Ett stort mönster - varavJag är en del - kanske min grejer rapade från någon bortglömd stjärna, som enär rapningar där. Eller se dem med större öga Palomar, rusar allabortsett från vissa gemensam utgångspunkt när de var kanske alla tillsammans.Vad är mönstret, eller innebörden, eller * varför? * Det gör inte skadamysterium att veta lite om det. För mycket mer underbart är sanningen ännågra artister från det förflutna trott! Varför poeterna i föreliggande inte talaav det? Vilka män är poeter som kan tala om Jupiter om han var som en människa, menom han är en enorm snurrande sfär av metan och ammoniak måste vara tyst?
		-- Richard P. Feynman (1918-1988)

%
Om du tillåter dig själv att läsa betydelser i (snarare än dra betydelser utav) bevis kan du dra någon slutsats du vill.
		-- Michael Keith, "The Bar-Code Beast", The Skeptical Enquirer Vol 12 No 4 p 416

%
"Pseudokod kan användas i viss utsträckning för att underlätta upprätthållandetbehandla. Men pseudokod som är mycket detaljerad -närmar detaljnivån i koden själv - är inte avmycket användning som underhållsdokumentation. sådan detaljeraddokumentation måste upprätthållas nästan lika mycket som den kod,alltså en fördubbling av försörjningsbördan. Vidare, eftersom en sådanomfattande pseudokod är alltför störande att hållas inotering själv, måste det hållas i en separat mapp. Deresultat: Eftersom pseudokod - till skillnad från riktiga kod - behöver inte varabibehålls, kommer ingen att upprätthålla den. Det kommer snart att bli avdatum och alla kommer att ignorera det. (En gång gjorde jag en informellundersökning av 42 butiker som används pseudokod. Av dessa 42, 0 [noll!]fann att det hade något värde som underhållsdokumentation. "         --Meilir Sida-Jones, "The praktisk guide till Structured           Design ", Yourdon Press (c) 1988
		-- Michael Keith, "The Bar-Code Beast", The Skeptical Enquirer Vol 12 No 4 p 416

%
"Endast en hjärnskadade operativsystem skulle stödja uppgift växling och integöra enkla nästa steg att stödja multitasking. "
		-- George McFry

%
Sigmund Freud påstås ha sagt att i sista hand hela fältetpsykologi kan minska biologisk elektrokemi.
		-- George McFry

%
Trollkarlen sitter i sin barnstol och ser på världen med fördel.Han är på höjden av sin makt. Om han sluter ögonen, orsakar han världenatt försvinna. Om han öppnar ögonen, orsakar han världen att komma tillbaka. Omdet finns harmoni i honom, världen är harmonisk. Om rage splittrar hansinre harmoni, är enheten i världen krossade. Om önskan uppstår inomhonom, yttrar han magiska stavelser som orsakar det önskade objektet visas.Hans önskemål, hans tankar, hans gester, hans ljud kommandot universum.
		-- Selma Fraiberg, _The Magic Years_, pg. 107

%
Ett djur som vet vem det är, en som har en känsla av sin egen identitet, ären missnöjd varelse, dömd att skapa nya problem för sig själv förvaraktigheten av hans vistelse på den här planeten. Eftersom varken mus eller schimpansenvet vad som, han skonas alla besvärliga problem som följer dettaupptäckt. Men så snart det mänskliga djuret som frågade sig denna frågadykt upp, kastade han sig själv och sina ättlingar till en evighet av tviveloch grubblande, spekulation och sanningssökande som har eggade honom genomårhundraden som obevekligt som hunger eller sexuell längtan. Schimpansen som görinte vet att han existerar inte drivs för att upptäcka sitt ursprung och skonasden tragiska nödvändigheten av överväger sin egen ände. Och även om djuretpraktiker lyckas lära en schimpans att räkna hundra bananer elleratt spela schack, kommer schimpansen utveckla ingen vetenskap och han kommer att uppvisa någonuppskattning av skönhet, för den största delen av mänsklig visdom kan spårastillbaka till de eviga frågorna om början och slut, att strävan att gevilket innebär att hans existens, till livet självt.
		-- Selma Fraiberg, _The Magic Years_, pg. 193

%
En kommentar om tidtabeller: Ok, hur lång tid tar det?   För varje engagerad i första möten manager lägga en månad.   För varje chef som säger "analys dataflödet" lägga ytterligare en månad.   För varje unik slutanvändaren typ lägga en månad.   För varje okänt mjukvarupaket som skall användas lägga till två månader.   För varje okänd hårdvaruenhet lägga till två månader.   För varje 100 miles mellan utvecklare och installation lägga en månad.   För varje typ av kommunikationskanal lägga en månad.   Om en IBM stordator butik är inblandade och du arbetar på en icke-IBM      Systemet lägger 6 månader.   Om en IBM stordator butik är inblandade och du arbetar på en IBM      Systemet lägger 9 månader.Runda upp till närmaste halvåret.--Brad ShermanFörresten, är alla mjukvaruprojekt görs av iterativ prototyping.Vissa företag kallar sina prototyper "utsläpp", det är allt.
		-- Selma Fraiberg, _The Magic Years_, pg. 193

%
    UNIX Shell är det bästa fjärde generationens programmeringsspråk    Det är den UNIX-skal som gör det möjligt att göra program i en liten    fraktion av koden och tiden det tar i tredje generationens språk. I    skalet du bearbetar hela filer på en gång, i stället för bara en linje på en    tid. Och är en kodrad i UNIX skalet ett eller flera program,    som gör mer än sidor med instruktioner i en 3GL. Ansökan kan vara    utvecklats i timmar och dagar, snarare än månader och år med traditionell    system. De flesta av de andra 4GLs finns idag ser mer ut COBOL eller    RPG, den mest tråkiga av tredje generationens språk."UNIX Relational Database Management: Application Development i UNIX Miljö "av Rod Manis, Evan Schaffer, och Robert Jörgensen. Prentice Hall Software Series. Brian Kerrighan, rådgivare. 1988.
		-- Selma Fraiberg, _The Magic Years_, pg. 193

%
"Skratta när du kan, apa-boy."
		-- Dr. Emilio Lizardo

%
"Spöstraff kommer att fortsätta tills moral förbättras."
		-- anonymous flyer being distributed at Exxon USA

%
"Hej Ivan, kontrollera din sex."- Sidewinder missil jacka lapp, som visar en Sidewinder driver upp svansen av en rysk Su-27
		-- anonymous flyer being distributed at Exxon USA

%
"Fria marknader väljer för att vinna lösningar."
		-- Eric S. Raymond

%
"Jag ogillar företag som har en vi-är-the-high-präster-of-hårdvaru så you'll-like-vad-vi-ge-du attityd. Jag gillar råvarumarknaderna där järn-och-kisel gatuförsäljare vet att de existerar för att ge snabba leksaker för programtyperatt jag ska spela med ... "
		-- Eric S. Raymond

%
"Lust att förstöra är också en kreativ lust."- Bakunin[Ed. Observera - Jag skulle säga: Driften att förstöra kan ibland vara en kreativ lust].
		-- Eric S. Raymond

%
"En kommersiell, och i vissa avseenden en social, tvivel har inletts inom senaste året eller två, om det är rätt att diskutera så öppet säkerheten eller osäkerhet av lås. Många välmenande personer anta att diskus- sionen respekterar medel för förbryllande den förmodade säkerhet lås har en premie för oärlighet, genom att visa andra hur man vara oärlig. Detta är en i träda Lacy. Rogues är mycket angelägna i sitt yrke, och redan vet mycket mer än vi kan lära dem att respektera sina olika typer av skurkaktighet. skälmar visste en hel del om lockpicking långt innan låssmeder diskuterade det bland dem- själva, eftersom de har nyligen gjort. Om ett lås - låt det ha skett i vad- någonsin land, eller av vad Maker - är inte så okränkbar eftersom den har hittills bedömts vara, det är säkert av intresse för * ärliga * personer att veta detta faktum, eftersom * oärlig * är tämligen säker på att vara den första som tillämpa kunskapen i praktiken; och spridning av kunskap är nödvändig för att ge rent spel för dem som kan drabbas av okunnighet. Det kan inte vara alltför öron nestly manade att en bekant med verkliga fakta kommer i slutändan vara bättre för alla parter. "- Charles Tomlinson s Rudimentary avhandling om konstruktion av lås,   offentliggöras omkring 1850
		-- Eric S. Raymond

%
 När det gäller att låsa fattandet, det kan knappast vara en sådan sak som oärlighet avsikt: uppfinnaren producerar ett lås som han ärligt tror kommer har sådana och sådana kvaliteter; och han förklarar sin tro till världen. Om andra skiljer sig från honom i yttrande om dessa kvaliteter, är det öppet till dem att säga så; och diskussionen, sanningsenligt genomförts, måste leda till offentliga fördel: diskussionen stimulerar nyfikenhet och nyfikenhet stimulerat lates uppfinning. Ingenting annat än en partiell och begränsad syn på frågan skulle kunna leda till uppfattningen att skada kan leda till: om det finns skador, kommer det att vara mycket mer än uppvägas av bra. "- Charles Tomlinson s Rudimentary avhandling om konstruktion av lås,   publiceras omkring 1850.
		-- Eric S. Raymond

%
"Inte vill tyckas, men för att vara det bästa."
		-- Aeschylus

%
"Undersökning säger ..."
		-- Richard Dawson, weenie, on "Family Feud"

%
"Paul Lynde att blockera ..."
		-- a contestant on "Hollywood Squares"

%
"Little else matters än att skriva bra kod."
		-- Karl Lehenbauer

%
Att skriva bra kod är en värdig utmaning, och en källa till civiliserade glädje.
		-- stolen and paraphrased from William Safire

%
"Stupidity, som dygd, är sin egen belöning"
		-- William E. Davidsen

%
"Om en dator inte direkt kan ta itu med alla RAM-minne du kan använda, det är bara en leksak."
		-- anonymous comp.sys.amiga posting, non-sequitir

%
"Never skratta åt levande drakar, Bilbo du dåre!" sade han till sig själv, och det bleven favorit talesätt av hans senare, och passerat in ett ordspråk. "Du är inte allsgenom detta äventyr ännu ", tillade han, och det var ganska sant också.
		-- Bilbo Baggins, "The Hobbit" by J. R. R. Tolkien, Chapter XII

%
"En smutsig sinne är en glädje för evigt."
		-- Randy Kunkee

%
"Du kan inte lära sju fot."- Frank Layton, Utah Jazz baskettränare, på frågan varför han hade rekryterat   en sju-fot hög bilmekaniker
		-- Randy Kunkee

%
"En bil är bara en stor väska på hjul."
		-- Johanna Reynolds

%
"Historien är ett verktyg som används av politiker för att rättfärdiga sina avsikter."
		-- Ted Koppel

%
"Gozer den gozerian: Som vederbörligen utsedd representant för staden,länet och staten New York, beställer jag härmed att upphöra med all övernaturligaktiviteter på en gång och gå direkt till ursprungsorten ellernärmaste parallell dimension, beroende på vilket som är närmast. "
		-- Ray (Dan Akyroyd, _Ghostbusters_

%
Man måste komma ihåg att det finns inget svårare att planera, mertveksam till framgång, inte heller farligare att hantera, än att skapa ennya systemet. För initiativtagaren har fiendskap alla som vill dra nytta avbevarandet av de gamla institutionerna och endast ljummet försvarare ide som skulle tjäna på de nya.
		-- Machiavelli

%
Gudlån mig senilitet att acceptera det jag inte kan förändra,Den frustration att försöka förändra saker jag kan inte påverka,och visdom att avgöra skillnaden.
		-- Machiavelli

%
Först som till tal. Det privilegium vilar på antagandet attDet finns ingen proposition så enhetligt erkänt att det inte kan varalagligen utmanade, ifråga och diskuteras. Det behöver inte vila påden ytterligare förutsättningen att det inte finns några påståenden som inte ärifrågasättas; det är tillräckligt, även om det finns, att i slutändan är detvärre att undertrycka oliktänkande än att riskera att kätteri. varför dethar om och om igen utan villkor proklamerade att det finnsinga gränser för förmånen såvitt ord försöker påverka endast åhörare "övertygelse och inte deras beteende. Problemet är detta beteende är nästanalltid baserade på någon tro, och att ändra åhöraren troi allmänhet i viss utsträckning ändra sitt beteende, och kan även framkallagenomföra att lagen förbjuder.[Jfr Lärt Hand, The Spirit of Liberty, University of Chicago Press, 1952;Konsten och Craft of döma: Besluten som domare Learned Hand,redigeras och kommenterad av Hershel Shanks, The MacMillian Company, 1968.]
		-- Machiavelli

%
Den sena upproret i Massachusetts har gett mer larm än vad jag tror detborde ha gjort. Räkna ut att en revolt i 13 stater under11 år, är men en för varje stat i ett och ett halvt sekel. inget landbör vara så länge utan en.
		-- Thomas Jefferson in letter to James Madison, 20 December 1787

%
"Nio år av balett, skitstövel."- Shelley Long, den onde efter att ha gjort ett hopp över en klyfta som han   kunde inte helt, i "Outrageous Fortune"
		-- Thomas Jefferson in letter to James Madison, 20 December 1787

%
Du är i en labyrint av UUCP anslutningar, alla lika.
		-- Thomas Jefferson in letter to James Madison, 20 December 1787

%
"Om den mannen i PTL är en sådan healer, varför kan han inte göra sin fru frisyr gå ner? "
		-- Robin Williams

%
8) Använd sunt förnuft i routing kabel. Undvik omslag koaxial runt källor     starka elektriska eller magnetiska fält. Linda inte kabeln runt     fluorescerande ljus förkopplingsdon eller cyklotroner, till exempel.- Ethernet Head produkt, information och installationshandbok,   Bell Technologies, sid. 11
		-- Robin Williams

%
"Vad ett konstigt är Usenet, sådan grossist produktion av gissningar frånen sådan obetydlig investering i själva verket. "
		-- Carl S. Gutekunst

%
VMS måste dö!
		-- Carl S. Gutekunst

%
MS-DOS måste dö!
		-- Carl S. Gutekunst

%
OS / 2 måste dö!
		-- Carl S. Gutekunst

%
Pournelle måste dö!
		-- Carl S. Gutekunst

%
Garbage in, Gospel ut
		-- Carl S. Gutekunst

%
"Att mot tortyr borde vara en slags multipartisan sak."
		-- Karl Lehenbauer, as amended by Jeff Daiell, a Libertarian

%
"Fakta är dumma saker."- President Ronald Reagan   (En blooper från sitt tal vid '88 GOP-konventionen)
		-- Karl Lehenbauer, as amended by Jeff Daiell, a Libertarian

%
"Argumentet att den bokstavliga historien om Genesis kan kvalificera som vetenskapkollapsar på tre viktiga skäl: kreationisternas behov av att åberopamirakel för att komprimera händelserna i jordens historia iden bibliska loppet av några tusen år; deras ovilja attöverge fordringar klart motbevisas inklusive påståendet att allafossil är produkter av Noas flod; och deras tillit distorsion,misquote, halv-citat och citat ur sitt sammanhang för att karakteriseraidéer sina motståndare. "- Stephen Jay Gould, "The Bedömning på kreationism",   Den Skeptical Inquirer, vintern 87/88, sid. 186
		-- Karl Lehenbauer, as amended by Jeff Daiell, a Libertarian

%
"Ett uns av förebyggande är värt ett ton av kod."
		-- an anonymous programmer

%
"IBM" öppen "innebär att det finns ett minimum av interoperabilitet mellan några av derasutrustning."
		-- Harv Masterson

%
"Tänk på en dator som hårdvara du kan programmera."
		-- Nigel de la Tierre

%
"Om du äger en maskin, är du i sin tur ägs av det, och tillbringa din tid betjänar det ... "
		-- Marion Zimmer Bradley, _The Forbidden Tower_

%
"Allt bör göras så enkelt som möjligt, men inte enklare."
		-- Albert Einstein

%
"Kortläsare? Behöver vi inte några stinkande kortläsare."- Peter da Silva (vid National Academy of Sciences, 1965, i en   särskilt levande fantasi)
		-- Albert Einstein

%
Din goda natur kommer att ge obegränsad lycka.
		-- Albert Einstein

%
Semper Fi, dude.
		-- Albert Einstein

%
Spänning och fara väntar din induktion till spår plikt! Som ett spårämne,du måste befria datornät av slemmiga, kriminella data tjuvar.De är svåra och de åtgärder som blir tufft, så se upp! utnyttja alladina kunskaper kommer du antingen få din man eller du bli bränd!
		-- advertising for the computer game "Tracers"

%
"En hel broderskap bandnings Wall-Street-bundna ungdom Hell -. Dettakommer att bli ett blodbad! "
		-- Post Bros. Comics

%
"Grannar !! Vi fick grannar! Är vi inte tänkt att ha några grannar, ochJag var bara tvungen att skjuta en. "
		-- Post Bros. Comics

%
"Gotcha, snor halsade du weenies!"
		-- Post Bros. Comics

%
. SPÄCKA - vt, för att blanda; diversifiera
		-- Webster's New World Dictionary Of The American Language

%
"Alla talar om vädret men ingen gör något åt ​​det."
		-- Mark Twain

%
"Hur många Teamsters tar det att skruva i en glödlampa?"   "Femton !! Har du problem med det?"
		-- Mark Twain

%
"Om du inte var min lärare, skulle jag tror att du tagit bort alla mina filer."- En anonym UCB CS student, en lärare som hade skrivit "rm -i *" till   bli av med en fil med namnet "f" på ett Unix-system.
		-- Mark Twain

%
"De hetaste platserna i helvetet är reserverade för dem som, i tider av moraliskkris, bevarat sin neutralitet. "
		-- Dante

%
"Mediet är budskapet."
		-- Marshall McLuhan

%
"Mediet är massagen."
		-- Crazy Nigel

%
"Visa mig en god förlorare, och jag ska visa dig en förlorare."
		-- Vince Lombardi, football coach

%
"Det kan hjälpa om vi körde MBA av Washington."
		-- Admiral Grace Hopper

%
Uppdateras av en kort blackout, fick jag till mina fötter och gick bredvid.
		-- Martin Amis, _Money_

%
De fjädrande dörrar skildes och jag stapplade ut i lobbyn teak och flimmer.Uniformerade män stod oberört som vaktposter i deras dike. jag slogmin nyckel på skrivbordet och nickade allvarligt. Jag var lastad nog att vara oförmögen attberätta om de kunde berätta jag laddades. Skulle de tänka? Jag var verkligenalltför laddad till vård. Jag flyttade till dörren med boxy, schlep axlade framsteg.
		-- Martin Amis, _Money_

%
Jag ber bara en sak. Jag förstår. Jag är mogen. Och det är inte mycket attfråga. Jag vill komma tillbaka till London, och spåra henne, och vara ensam med minSelina - eller ens ensam, fan, bara nära henne, tillräckligt nära för attlukta hennes hud, för att se fläckiga bandet hennes lemony ögon, gjutningav sin konstfulla läppar. Bara för några dyrbara sekunder. Bara tillräckligt länge för attsätta i en bra, ren punch. Det är allt jag ber.
		-- Martin Amis, _Money_

%
"Love kan misslyckas, men artighet kommer previal."
		-- A Kurt Vonnegut fan

%
New York är en djungel, de berätta. Du kan gå vidare och säga attNew York är en djungel. New York * är en djungel. * Under kolumnernaden gamla regnskogen, gjord av smält makadam, medelvärdet Limpopo av översvämmasNinth Avenue bär en arg argosy av crocs och drakar, tiger fisk, bullermaskiner, svettningar regnmakare. På hörnen står witchdoctors ochheadhunters, porlande voodoo-män - de infödda, djungeln marta infödda.Och på natten, under ekvatorial överväxt och värmehållande molntäcka, hör du trasiga papegoja-hoot och monkeysqueak av sirener,och sedan skjuter blomma att avvärja monster. Noggrann: gatorna ärvuxit med gropar och nät och fällor. Hyra en guide. Packa ormbettGook och din blowdart serum. Ta det på allvar. Du måste få enbitars djungel-wise.
		-- Martin Amis, _Money_

%
Nu var jag på väg, i min varma bur, ned mot köttmarknaden land påspetsen av West Village. Här rött tegel lager dubbelt så kadavergallerier och råtta nässelfeber, Manhattan fauna som söker sin nödvändiganivå, levande eller död. Även här hittar du de tunga risknippe hangouts,Spike, Water Closet, Moder Load. Ingen vet vad som händerpå dessa platser. Endast de tunga fagots vet. Även Fielding verkar någotvag i frågan. Du får zapped och piskades och dumpas på - genomnästan någons standarder, har du verkligen fruktansvärd tid. Genomsnittetbeskyddare anländer till Spike i en taxi men behöver gå tillbaka till sin strumpaitu. Och sedan nästa natten han dyker upp mer. de schackelsig till ställningar, de hyllas i urinoarer. Deras föräldrar har en hel delförklarar att göra, om du vill ha min åsikt, särskilt mammor. Förlåtatt peka du damer ut så här men historien måste börja någonstans.En craving för hourly mord - det kan inte ville. Sålänge,Fielding säger, naturen ser på och knackar hennes fot och klicktungan. Alltid en förkämpe för monogami, hon kokar ihop några tjusiganya sjukdomar. Hon bara inte kommer att stå för det.
		-- Martin Amis, _Money_

%
"Du försökte det bara för en gångs skull, fann det okej för sparkar, men nu du ta reda på har du en vana som sticker, du är en orgasm missbrukare, du är alltid på det, och du är en orgasm missbrukare. "
		-- The Buzzcocks

%
"Det finns ingen distinkt amerikansk kriminell klass utom kongressen."
		-- Mark Twain

%
"Du betalar för att veta vad du verkligen tror."
		-- J. R. "Bob" Dobbs

%
"Vi lever i en mycket knasig tid."
		-- Herb Blashtfalt

%
"Slå blå dunster egna ögon!"
		-- J. R. "Bob" Dobbs

%
"Okej," Bobby sa, att få kläm på det, "vad är matrisen? Omhon är ett däck, och Danbala är ett program, vad är cyberrymden? "  "Världen", sa Lucas.
		-- William Gibson, _Count Zero_

%
"Våra repriser är bättre än deras."
		-- Nick at Nite

%
Livet är ett spel. Pengar är hur vi håller poäng.
		-- Ted Turner

%
"Betala ingen uppmärksamhet åt mannen bakom gardinen."
		-- The Wizard Of Oz

%
"Betala ingen uppmärksamhet åt mannen bakom gardinen."
		-- Karl, as he stepped behind the computer to reboot it, during a FAT

%
"Det är inte så mycket saker som vi inte vet att få oss i trubbel. Det ärsaker som vi vet att det är inte så. "
		-- Artemus Ward aka Charles Farrar Brown

%
"Inte rabatt flygande grisar innan du har bra luft försvar."
		-- jvh@clinet.FI

%
"I det långa loppet, blir varje program rokokor, och sedan spillror."
		-- Alan Perlis

%
"Pok POK pok, P'kok!"
		-- Superchicken

%
Levande fritt eller bor i Massachusetts.
		-- Superchicken

%
"Du kan inte få mycket långt i denna värld utan ditt underlag är det först."
		-- Arthur Miller

%
"Flyg Bokningssystem avgöra om du finns. Om informationenär inte i deras databas, då du helt enkelt inte får gå någonstans. "
		-- Arthur Miller

%
"Vad folk har reducerats till är endast 3-D representationer av sin egendata."
		-- Arthur Miller

%
"The Avis WIZARD avgör om du får köra bil. Ditt huvud kommer inte rörakudde av en Sheraton om datorn säger att det är okej. "
		-- Arthur Miller

%
"De vet ditt namn, adress, telefonnummer, kreditkortsnummer, vemär att köra bilen "för försäkring", ... din körkortsnummer. idelstaten Massachusetts, är detta samma nummer som används för socialaSäkerhet, om du motsätter sig sådan användning. I så fall är du tilldelas ennummer och du bor alltid mer på listan över "konstiga människor som inte gerut deras socialförsäkringsnummer i Massachusetts. "
		-- Arthur Miller

%
"Data är en mycket som människor: Det föds Matures gifter sig till andra uppgifter,..skild. Blir gamla. En sak som det inte gör är att dö. Det måste avlivas. "
		-- Arthur Miller

%
"Människor bör ha tillgång till de uppgifter som du har om dem. Det bör vara en process för dem att utmana eventuella felaktigheter. "
		-- Arthur Miller

%
"Även om polackerna lider officiell censur, en genomgripande hemlighetpolis och lagar liknande dem i Sovjetunionen, det finnstusentals jordiska publikationer, en juridisk oberoendeKyrka, privata jordbruk och östblocket första och endaoberoende facklig federation, NSZZ Solidarnosc, som ärett dotterbolag till både Internationella konfederationen för friaFackföreningar och World Confederation of Labor. Det finnsbokstavligen en värld av skillnad mellan Polen - även i sinnuvarande kollaps - och sovjetiska samhället på toppen avdess "glasnost." Denna skillnad har legat kvar på brakosta av polackerna sedan 1944.- David Phillips, SUNY på Buffalo, om upprättande av en   gateway från EARN (Eurpoean Academic Research Network)   till Polen
		-- Arthur Miller

%
"Det finns också en blomstrande oberoende studentrörelse iPolen och sålunda finns det en stark möjlighet (men ingengarantera) för att göra en earn-Polen länk, bör det någonsin kommaom en verklig länk - inte ett dammsugarmunstycke för enBloc informationsinsamling apparat ransone till förstapparatjiks. "- David Phillips, SUNY på Buffalo, om upprättande av en   gateway från EARN (Eurpoean Academic Research Network)   till Polen
		-- Arthur Miller

%
"Inte förlora dina kunskaper att människans rätt egendom är en upprätt hållning,en oförsonlig sinne, och ett steg som reser obegränsade vägar. "
		-- John Galt, in Ayn Rand's _Atlas Shrugged_

%
Inte panik.
		-- John Galt, in Ayn Rand's _Atlas Shrugged_

%
Felet slutar här.
		-- John Galt, in Ayn Rand's _Atlas Shrugged_

%
Felet börjar här.
		-- John Galt, in Ayn Rand's _Atlas Shrugged_

%
"Varför slösa negativ entropi på kommentarer, när du kan använda sammaentropi för att skapa fel i stället? "
		-- Steve Elias

%
"Den patologi är att vill ha kontroll, inte att du någonsin få det, på grund avNaturligtvis aldrig göra. "
		-- Gregory Bateson

%
"Din rumpa är min."
		-- Michael Jackson, Bad

%
Skicka den.
		-- Michael Jackson, Bad

%
"När de går upp, vem bryr sig när de kommer ner? Det är inte min avdelning."
		-- Werner von Braun

%
"När det enda verktyg man har är en hammare, tenderar man att behandla allt som omdet var en spik. "
		-- Abraham Maslow

%
"Imitation är den ärligaste formen av TV."
		-- The New Mighty Mouse

%
"Den mindre av två onda ting - är ond."
		-- Seymour (Sy) Leon

%
"Det är ingen svett, Henry. Russ gjort det tillbaka till Bugtown innan han dog. Så han skaregenerera i ett par dagar. Det är bara hemskt slarvigt av honom att bli dödad iförsta hand. Humph! "
		-- Ron Post, Post Brothers Comics

%
"En ärlig gud är den ädlaste människans verk. ... Gud har alltid liknade hanskreatörer. Han hatade och älskade vad de hatade och älskade och han var alltidfinns på sidan av makthavarna. ... De flesta av gudarna var nöjda medoffra, och lukten av oskyldigt blod har någonsin ansetts vara en gudomligparfym."
		-- Robert G. Ingersoll

%
"Vi är inte försöker kedjan framtiden, men att frigöra den nuvarande. ... Vi ärförespråkare undersöknings, utredning, och tanke. ... Det är stors att tänkaoch undersöka själv än att upprepa en trosbekännelse. ... Jag ser för dagennär * anledning *, throned på världens hjärnor ska vara kungen av Kings ochGud Gods.
		-- Robert G. Ingersoll

%
"Jag tror verkligen att läran om helvetet föddes i de glittrande ögonenav ormar som körs i fruktansvärda spolar tittar på sina byten. Jag trordet föddes med yelping, tjutande, morrande och morrande av vilda djur ...Jag föraktar det, jag trotsar det, och jag hatar det. "
		-- Robert G. Ingersoll

%
"Är detta förspel?"   "Nej, det är Nuke Strike. Förspel har usel grafik. Slå mig igen."
		-- Duckert, in "Bad Rubber," Albedo #0 (comics)

%
egrep mönster är fulla reguljära uttryck; den använder en snabb deterministiskalgoritm som ibland behöver exponentiell utrymme.
		-- unix manuals

%
"Ett sinne är en fruktansvärd sak att ha läcker ut öronen."
		-- The League of Sadistic Telepaths

%
"Livet suger, men det är bättre än alternativet."
		-- Peter da Silva

%
Om detta är en tjänsteekonomi, varför är tjänsten så illa?
		-- Peter da Silva

%
"Jag förväntar mig en kemisk bot för psykopat beteende från 10:00 i morgon,eller jag har dina tarmar för spaghetti. "
		-- a comic panel by Cotham

%
"Även om du är på rätt spår, du får köra över om du bara sitter där."
		-- Will Rogers

%
"Ett öppet sinne har men en nackdel: det samlar smuts."
		-- a saying at RPI

%
"Geeksna ärva jorden."
		-- Karl Lehenbauer

%
"Akta dig för programmerare som bär skruvmejslar."
		-- Chip Salzenberg

%
"Elvis är min copilot."
		-- Cal Keegan

%
"Den grundläggande principen för vetenskap, definitionen nästan, är detta:enda test av giltigheten av någon aning är experiment. "
		-- Richard P. Feynman

%
Hur många Unix hacka tar det att byta en glödlampa?   Låt oss se, kan du använda ett skalskript för det eller behöver det ett C-program?
		-- Richard P. Feynman

%
"Hata inte mig eftersom jag är vacker. Hatar mig för att jag är vacker, smartoch rik. "
		-- Calvin Keegan

%
"Hela problemet med världen är att dårar och fanatiker är alltid såvissa av sig själva, men klokare människor så fulla av tvivel. "
		-- Bertrand Russell

%
ser alltid över axeln eftersom alla tittar på och plottamot dig.
		-- Bertrand Russell

%
"Låt oss fördöma till hellfire alla dem som inte håller med oss."
		-- militant religionists everywhere

%
Bäbis ombord.
		-- militant religionists everywhere

%
"Nettoresultatet är ett system som inte bara är binärt kompatibla med 4,3 BSD,men är även bug för kryp kompatibla i nästan alla funktioner. "- Avadit Tevanian, Jr., "Arkitektur-oberoende virtuella minneshantering   Parallell och distribuerade miljöer: Mach Approach "
		-- militant religionists everywhere

%
"Antalet Unix installationer har vuxit till 10, med mer väntat."
		-- The Unix Programmer's Manual, 2nd Edition, June, 1972

%
"Engineering utan management är konst."
		-- Jeff Johnson

%
"Jag är inte en gud, jag var felciterad."
		-- Lister, Red Dwarf

%
Hjärna off-line, var god vänta.
		-- Lister, Red Dwarf

%
-! - UUNet socker karl | "Vi har följt dina framsteg med betydande- Karl@sugar.uu.net | intresse, att inte säga förakt "-. Zaphod Beeblebrox IV- Usenet BBS (713) 438-5018th-th-th-th-det är allt, folks!----------- Skära här, glöm inte att beröva skräp i slutet, alltför -------------"Psyko ?? Jag trodde att detta var en naken rap session !!!"
		-- Zippy

%
Har du roligt ännu?
		-- Zippy

%
"De allra flesta framgångsrika stora brott mot egendombegås av individer som missbrukar förtroendeuppdrag. "
		-- Lawrence Dalzell

%
"Kanske jag piskning ett sugrör sill i mitten av strömmen, men mot bakgrund avvad som är känt om den gränslösa säkerhetsproblem, verkar det kraftigtför farligt för universitets folk att köra med huvudet i sanden. "
		-- Peter G. Neumann, RISKS moderator, about the Internet virus

%
"Seed mig, Seymour"
		-- a random number generator meets the big green mother from outer space

%
"Köp mark. De har slutat göra det."
		-- Mark Twain

%
"Öppna pod bay dörrar, HAL."
		-- Dave Bowman, 2001

%
"Det var ingen skillnad mellan beteendet hos en gud och verksamhetren slump ... "
		-- Thomas Pynchon, _Gravity's Rainbow_

%
... Saure verkligen visar sig vara en skicklig på den svåra konsten att papryomancy,förmågan att sia genom överväger hur människor rulla kylfartyg -formen, slickande mönster, rynkor och veck eller frånvaro däravi tidningen. "Du kommer snart att vara kär" sez Saure, "se, denna linje här.""Det är lång, är inte den gör att medelvärdet -?" "Längd är oftast intensitet.Inte tid. "
		-- Thomas Pynchon, _Gravity's Rainbow_

%
Gå vidare, kapitalisera T på teknik, avguda det om det får dig att kännamindre ansvariga - men det sätter du in med kastrerad, bror, in medeunucker hålla harem av vår stulna Earth för stel och glädjelöshardons mänskliga sultaner, för människors elit utan rätt alls vara där deär - "
		-- Thomas Pynchon, _Gravity's Rainbow_

%
... Den rådande katolska lukt - rökelse, vax, århundraden av mild bräkandefrån läppar flocken.
		-- Thomas Pynchon, _Gravity's Rainbow_

%
... På den tiden [1960], projicerade Bell Laboratories forskare somdatorhastigheter så höga som 30 miljoner flyttalsberäkningar perandra (megaflops) skulle behövas för arméns ballistiska missilerförsvarssystem. Många dataexperter - inklusive en National AcademyVetenskapsakademien panel - sade uppnå dessa hastigheter, även med hjälp av multipelprocessorer, var omöjligt. Idag, den nya generationens superdatorer fungerarvid miljarder operationer per sekund (gigaflop).
		-- Aviation Week & Space Technology, May 9, 1988, "Washington Roundup", pg 13

%
säkerhetskopiering: alltid i säsong, aldrig omodernt.
		-- Aviation Week & Space Technology, May 9, 1988, "Washington Roundup", pg 13

%
"Det fanns en vag, obehaglig manginess om hans utseende, han på något sättverkade smutsiga, men en nära blick visade honom så noggrant rakat som enskådespelare, och klädd i oklanderlig linne. "
		-- H. L. Mencken, on the death of William Jennings Bryan

%
Arbetet var omöjligt. Nördar hade brutit min ande. De hade gjort förmånga saker som är fel. Det var aldrig så här för Mencken. Han levde somen preussisk spelare - svettningar värre än Bryan på vissa nätter och fullareän Judas på andra. Det var allt en dehumanized mardröm ... och dessaraddled cretins har mage att klaga mina deadlines.
		-- Hunter Thompson, "Bad Nerves in Fat City", _Generation of Swine_

%
"Denna generation kan vara en som kommer att möta Armageddon."
		-- Ronald Reagan, "People" magazine, December 26, 1985

%
... Kabeln hade klarat oss; skålen var det enda hoppet, och så småningomVi var alla tvungna att vända sig till den. Vid sommaren av '85, hade dalen merparabolantenner per capita än en eskimå by på norra sluttningen avAlaska.Gruvan var en av de sista att gå i. Jag hade varit nervös redan från början omriskerna med alltför mycket input, vilket är ett mycket verkligt problem med dessasaker. Titta på TV blir en heltidsarbete när du kan skanna 200 kanalerhela dagen och hela natten och fortfarande har möjlighet att stansa Night Dreamsi video maskin, om resten av världen verkar tråkigt.
		-- Hunter Thompson, "Full-time scrambling", _Generation of Swine_

%
"Ring omedelbart. Tiden rinner ut. Vi båda behöver göra någotmonstruösa innan vi dör. "
		-- Message from Ralph Steadman to Hunter Thompson

%
"Det enda sättet för en reporter att titta på en politiker är nere."
		-- H. L. Mencken

%
"Du behöver inte gå ut och sparka en galen hund. Om du har en galen hund med rabies, duta en pistol och skjuta honom. "
		-- Pat Robertson, TV Evangelist, about Muammar Kadhafy

%
David Brinkley: Den dagliga astrologiska diagram är just där, i min  dom, de tillhör, och det är på den komiska sidan.George Will: Jag tror inte att astrologi hör även på komiska sidor.  De serier gör ingen sanning anspråk.Brinkley: Var skulle du säga?Kommer: Jag skulle inte sätta det i tidningen. Jag tror att det är transparent skräp.  Det är en återspegling av en idé som vi ut från det västerländska tänkandet i  sextonde århundradet, att vi är i mitten av en omtänksam universum. Vi är  inte i mitten av universum, och det bryr sig inte. Stjärnans anpassning  vid tiden för vår födelse - det är struntprat. Det är inte roligt att  har det inkräktat bland människor som har kärnvapen.Sam Donaldson: Detta är inte något nytt. Guvernör Ronald Reagan svors  strax efter midnatt i sin första sikt i Sacramento, eftersom stjärnorna  sa att det var ett gynnsamt tid.Will: De [horoskop] är fullkomlig laga banaliteter. De kan gälla  vem som helst och vad som helst.Brinkley: När är den exakta tidpunkten [födelse]? Jag tror inte att sjuksköterskan är  står där med ett stoppur och ett anteckningsblock.Donaldson: Om vi ​​fattar beslut baserat på stjärnorna - det är en cockamamie  sak. Folk vill veta.- "Denna vecka" med David Brinkley, ABC Television, Söndag 8 maj, 1988,   utdrag ur en diskussion om astrologi och Reagan
		-- Pat Robertson, TV Evangelist, about Muammar Kadhafy

%
Det rapporterade gripa astrologi i Vita huset har orsakat mycketmunterhet. Det är inte roligt. Astro rotvälska, vilket innebär astrologii allmänhet, har ingen plats i en tidning, att inte tala om regeringen. Till skillnad från serier,som är en del av en tidningens ofarlig nöje och gör inga sanningsanspråk,astrologi är ett bedrägeri. Tanken att det blir en utfrågning i regeringen ärförfärande.
		-- George Will, Washing Post Writers Group

%
Astrologi är den skir hokum. Denna pseudovetenskap har funnits sedandagen kaldéerna och babylonierna. Det är lika falsk som numerologi,phrenology, palmistry, alkemi, läsningen av teblad, och praktikspådom av inälvorna på en get. Ingen seriös person kommer att köpauppfattningen att våra liv påverkas individuellt genom förflyttning avavlägsna planeter. Detta är sågspån blarney av karnevalen halvvägs.
		-- James J. Kilpatrick, Universal Press Syndicate

%
En seriös offentlig debatt om giltigheten av astrologi? En allvarlig troendei Vita huset? Två av dem? Ge mig en paus. Vad kvävs min skrattär att bilden passar. Reagan har alltid uppvisat en fey likgiltighet motvetenskap. Fakta, samma siffror, rulla ut ryggen. Och vi har alla kommit tillacceptera den. Denna gång var stjärnorna som blev en allvarlig fråga .... Inteså länge sedan var det Reagans stöd av kreation .... Creationists faktisktfick samma tid med evolutionister. Allmänheten skulle vara öppentill anspråk paleontologer och fundamentalister, som om de två varvetenskapliga kollegor .... Det har stått klart länge att presidentenär främmande för vetenskapen ... I allmänhet är dessa attityder faller på vänlig amerikansktorv .... Men vid ytterkanterna, denna skepsis om vetenskap lätt vändertill ett slags naiv godkännande av nonscience, eller till och med nonsens. Det sammamänniskor som tvivlar experter kan också tro alla kvacksalveri, från fördelarna medLaetrile mot öga av newt till förflyttning av planeter. Vi förlorar förmågan attgöra rationella - vetenskapliga - domar. Det är i alla fall.- Ellen Goodman, The Boston Globe tidningen företaget Washington Post Writers    Grupp
		-- James J. Kilpatrick, Universal Press Syndicate

%
Skådespelet av astrologi i Vita huset - det styrande centrumvärldens största vetenskapliga och militära makt - är så skrämmande attdet trotsar förståelse och ger skäl för stor förskräckelse. Det lättastesvaret är att skratta bort det, och att hänge sig åt wisecracks om CivilTjänste betyg för horoskop beslutsfattare och palm läsare och om Reaganfrågade Michail Gorbatjov för hans tecken. En smittsam gott mod ärkännetecknande för detta ordförandeskap, även när det gäller de mest dystra frågor.Men den här gången, är det inte roligt. Det är vanligt skrämmande.- Daniel S. Greenberg, redaktör, _Science och regerings Report_, skriver i   "Newsday", 5 maj 1988
		-- James J. Kilpatrick, Universal Press Syndicate

%
[Astrologi är] 100 procent hokum, Ted. I själva verket, den första upplaganav Encyclopaedia Britannica, skriven i 1771 - 1771! - Sade att dettatrossystem är ett ämne för länge sedan förlöjligad och avskydda. Vi har att göra medövertygelser som går tillbaka till de gamla babylonierna. Det finns inget där ....Det låter väldigt lik vetenskap, det låter som astronomi. Det har fått tekniskvillkor. Det har fått jargong. Det förvirrar allmänheten .... Astrologen är ganskaglib, förvirrar allmänheten använder termer som kommer från vetenskapen, kommer frånmetafysik, kommer från en mängd olika områden, men de betyder egentligen ingenting. DeFaktum är att astrologiska föreställningar gå tillbaka åtminstone 2500 år. Nu närbör vara en tillräckligt lång tid för astrologer att bevisa sin sak. Dehar inte visat sig vara fallet .... Det är helt enkelt rappakalja. Faktum är, att det finnsingen teori för det, det finns inga observationsdata för det. Det har testatsoch testas under århundraden. Ingen har någonsin hittat någon giltighet till den påalla. Det är inte ens nära till en vetenskap. En vetenskap måste vara repeterbart, detmåste ha en logisk grund, och det måste vara potentiellt sårbara -du testa det. Och i att astrologi är verkligen något helt annat.- Astronomen Richard Berendzen, VD, American University, på ABC    Nyheter "Night" 3 maj 1988
		-- James J. Kilpatrick, Universal Press Syndicate

%
Med nyheten att Nancy Reagan har hänvisat till en astrolog vid planeringmakens schema, och rapporter om kalifornier evakuerings Los Angelespå styrkan av en förutsägelse från en sextonde-talet läkare ochastrolog Michel de Notredame, bilden av den amerikanska som en vetenskaplig ochteknisk nation har tagit lite av en misshandel på sistone. Tyvärr, såhappenings kan inte avfärdas som hugskott. De är manifestationerav en väletablerad "anti-science" tendensen i USA som i slutändan,kan hota landets ställning som en teknologisk makt. . . . Demanifestera utbredd önskan att avvisa rationalitet och ersätta en serieav quasirandom tro för att förstå universum bådar intebra för en nation djupt oroad över sin förmåga att konkurrera med sinindustriella jämlikar. Till den grad att den återspeglar tänker på enbetydande del av allmänheten, denna synpunkt uppmuntrar okunnighetoch, faktiskt, förakt för vetenskap och rationella metoder att närma sigsanning. . . . Det blir uppenbart att om USA inte plocka upp sigsnart och ägna vissa ansträngningar att utbilda unga effektivt sin förhoppning omupprätthålla ett sken av ledarskap i världen kan vila, paradoxalt nog,med en ny våg av tekniskt intresserade och utbildade invandrare som intelider av anti-vetenskap sjukdom frodas i en till synes ruttnande samhälle.
		-- Physicist Tony Feinberg, in "New Scientist," May 19, 1988

%
mirakel: ett extremt utestående eller ovanlig händelse, ting, eller prestation.
		-- Webster's Dictionary

%
"Den programmerare är en skapare av universum som han ensam är ansvarig. Universum av praktiskt taget obegränsad komplexitet kan vara skapas i form av datorprogram. "
		-- Joseph Weizenbaum, _Computer Power and Human Reason_

%
"Om koden och kommentarerna håller, då båda är antagligen fel."
		-- Norm Schryer

%
"Må din framtid endast begränsas av dina drömmar."
		-- Christa McAuliffe

%
"Det är bättre för civilisationen att gå ner i avloppet än att varakommer upp det. "
		-- Henry Allen

%
"Livet börjar när du kan tillbringa fritiden programmering i stället förtittar på TV."
		-- Cal Keegan

%
"Vi gör aldrig påståenden, fröken Taggart", säger Hugh Akston. "Det ärden moraliska brott utmärkande för våra fiender. Vi berättar inte - vi * Visa *.Vi hävdar inte - vi * bevisa * ".
		-- Ayn Rand, _Atlas Shrugged_

%
"Jag minns när jag var liten brukade jag komma hem från söndagsskolan och min mamma skulle bli full och försöka göra pannkakor. "
		-- George Carlin

%
"Min far? Min far lämnade när jag var ganska ung. Jo faktiskt, han ombads att lämna. Han hade svårt metaboliserar alkohol. "
		-- George Carlin

%
"Jag slår på TV: n. Jag ser en ung kvinna som går under täckmantelför att vara en kristen, känd över hela landet, klädd i huden tätaskinnbyxor, skakningar och vickar hennes höfter i takt och rytmmusik som strobe lampor slår sina mönster över scenen ochbandet spelar den samtida rocksound som inte kan skiljas frånlåtar från Grateful Dead, Beatles, eller någon annan. Och du kan provaatt berätta detta är av Gud och att det leder människor till Kristus, men jagvet bättre.- Jimmy Swaggart, hycklande sexuell pervers och TV predikant, beskriver sig själv pornografi missbrukare, "Två synvinklar." Christian "rock and roll", Evangelisten, 17 (8): 49-50.
		-- George Carlin

%
"Så kallade kristen rock.... Är en djävulsk kraft underminera kristendom inifrån."- Jimmy Swaggart, hycklare och TV predikant, beskriver sig själv som pornografi missbrukare, "Två synvinklar:." Christian "rock and roll", evangelisten, 17 (8): 49-50.
		-- George Carlin

%
"Någon försöker generera slumptal med deterministiska sätt är,Naturligtvis lever i ett tillstånd av synd. "
		-- John Von Neumann

%
"Du måste ha en IQ på minst en halv miljon." - Popeye
		-- John Von Neumann

%
"Frihet är fortfarande den mest radikala idén om alla."
		-- Nathaniel Branden

%
Är du inte glad att du inte få alla regeringen du betalar för nu?
		-- Nathaniel Branden

%
"Jag lät aldrig min skolgång komma i vägen för min utbildning."
		-- Mark Twain

%
Dessa screamingly lustiga Gogs säkerställa ägare av X Ray Gogs att vara livetav någon part.
		-- X-Ray Gogs Instructions

%
En elev frågade befälhavaren om hjälp ... gör detta program körs frånArbetsbänk? Befälhavaren tog musen och pekade på en ikon. "Vad ärdetta? "frågade han. Studenten svarade" Det är musen ". Befälhavaren pressadekontroll Amiga-Amiga och träffade student på huvudet med Amiga ROM KernelManuell.
		-- Amiga Zen Master Peter da Silva

%
"Tack och lov för startups, utan dem vi aldrig skulle ha några framsteg."
		-- Seymour Cray

%
"Ut ur registret utrymme (ugh)"
		-- vi

%
"Dess brister trots, det finns mycket att säga till förmånjournalistik i det genom att ge oss yttrandet från outbildade,det håller oss i kontakt med okunskap i samhället. "
		-- Oscar Wilde

%
"Ada är PL / I försöker vara Smalltalk.
		-- Codoso diBlini

%
"De största hoten mot frihet lurar i smygande intrång av män av iver,välmenande men utan att förstå. "
		-- Justice Louis O. Brandeis (Olmstead vs. United States)

%
" 'Tis sant,' tis synd, och synd" tis "tis sant."- Poloniouius i Willie Shake s _Hamlet, Prince of Darkness_
		-- Justice Louis O. Brandeis (Olmstead vs. United States)

%
"Alla människor är så lycklig nu, deras huvuden grottkrypning. Jag är glad att deär en snögubbe med skyddande gummi hud "
		-- They Might Be Giants

%
"Obeslutsamhet är grunden för flexibilitet"
		-- button at a Science Fiction convention.

%
"Ibland vansinne är det enda alternativet"
		-- button at a Science Fiction convention.

%
"Ålderdom och förräderi kommer att slå ungdom och skicklighet varje gång."
		-- a coffee cup

%
"Det viktigaste i en människa är inte vad han vet, men vad han är."
		-- Narciso Yepes

%
"Allt vi får är möjligheter - att göra oss en eller annan sak."
		-- Ortega y Gasset

%
"Vi kommer att bli bättre och modigare om vi engagerar och fråga än om vi ägna sig åttomgångs infall som vi redan vet - eller att det är till någon nytta att försökavet vad vi inte vet. "
		-- Plato

%
"Att genomföra ett projekt, som ordets härledning antyder innebär att kasta enidé ut framför sig så att det får autonomi och uppfylls inte baraav de ansträngningar som dess upphovsman, men faktiskt, oberoende av honom också.
		-- Czeslaw Milosz

%
"Vi kan inte skjuta upp levande tills vi är redo. Den mest framträdande egenskaplivet är dess coerciveness; det är alltid angeläget, "här och nu", utan någoneventuell senareläggning. Livet avfyras på oss peka tomt. "
		-- Ortega y Gasset

%
"Därifrån till här, härifrån till dit, roliga saker finns överallt."
		-- Dr. Seuss

%
"När det gäller ödmjukhet, jag är den största."- Bullwinkle Moose
		-- Dr. Seuss

%
Kom ihåg att en int är inte alltid 16 bitar. Jag är inte säker, men om 80386 är ensteg närmare Intels slugfest med CPU kurva som är asymptotisktnärmar sig en riktig maskin, kanske en int har genomförts som 32 bitar avvissa Unix leverantörer ...?
		-- Derek Terveer

%
"I den mån jag kan höras av något, som kanske eller kanske inte bryr sigvad jag säger, frågar jag, om det är viktigt att du bli förlåten för någotdu kan ha gjort eller underlåtit att göra som kräver förlåtelse.Omvänt, om inte förlåtelse, men något annat kan krävas för attförsäkra alla möjliga nytta som du kan vara berättigad efterförstörelse av kroppen, ber jag att detta vad det nu kan vara,beviljas eller undanhålls, i förekommande fall kan vara, på ett sådant sätt attförsäkra din mottagning av nämnda förmån. Jag frågar detta i min egenskap avdin valda mellanhand mellan dig själv och det som inte kan varasjälv, men som kan ha ett intresse i fråga om dinmottagning så mycket som det är möjligt för dig att få av dettasak, och som kan på något sätt påverkas av denna ceremoni. Amen."Madrak i _Creatures av ljus och Darkness_, av Roger Zelazny
		-- Derek Terveer

%
"En akademisk spekulerade om en badande är vackerom det inte finns någon i skogen för att beundra henne. han gömdei buskarna för att ta reda på, som behäftat hans premissmen gjorde honom lycklig.Moral: Empirism är roligare än spekulationer ".
		-- Sam Weber

%
1 1 var en kapplöpningshäst, 2 2 var en 2. När en 1 1 1 ras, 2 2 1 1 2.
		-- Sam Weber

%
"Jag tänkte att det var denna förintelse, höger, och de enda kvar i livet var Donna Reed, Ozzie och Harriet, och Cleavers. "- Wil Wheaton förklarar varför alla i "Star Trek: The Next Generation"    är så trevligt
		-- Sam Weber

%
"Engineering möter konst på parkeringen och saker explodera."
		-- Garry Peterson, about Survival Research Labs

%
"Varför kan inte vi någonsin försöka lösa ett problem i det här landet utanen "War" på det? "- Rich Thomson, talk.politics.misc
		-- Garry Peterson, about Survival Research Labs

%
      ... Och innan jag visste vad jag gjorde, hade jag sparkade      skrivmaskin och kastade den runt i rummet och gjorde det tigga      barmhärtighet. Vid denna punkt skrivmaskin bad för mig att klä      honom i feminina kläder utan jag tryckte hans marginal frigivning      om och om igen tills skrivmaskin förlorade medvetandet.      För närvarande återfick jag medvetandet och insåg med skam vad      Jag hade gjort. Min skam är borta och nu är jag letar efter en      undergiven skrivmaskin, vilken färg som helst, eller modell. ingen elektrisk      skrivmaskiner tack!
		-- Rick Kleiner

%
Professionell brottning: balett för den vanliga människan.
		-- Rick Kleiner

%
"En idealist är en person som på märker att en ros luktar bättre än enkål, drar slutsatsen att det också kommer att göra bättre soppa. "- H.L. Mencken
		-- Rick Kleiner

%
   "Är dessa cocktail-servitrisen fingertecken?" Jag frågade Colletti som hanvisade oss dessa repor på bröstet. "Nej, de är på min rygg," Collettibesvaras. "Det är där ett fall av cocktail räkor föll på mig. Jag berättade för henneatt sakta ner lite, men du vet cocktail servitriser, de verkar haett sinne för sin egen. "- Den otroligt Monstrous, Mind-Rostning Summer of O.C. och Stiggs   National Lampoon, oktober 1982
		-- Rick Kleiner

%
"Ge aldrig i. Ge aldrig i. Aldrig. Aldrig. Aldrig."
		-- Winston Churchill

%
"Aldrig skriver malice det som orsakas av girighet och okunnighet."
		-- Cal Keegan

%
"Trots sin suffix, är skepticism inte en" ism "i betydelsen av en troeller dogma. Det är helt enkelt ett sätt att angripa problemet för att tala om vad som ärförfalskade och vad som är äkta. Och en erkännande av hur dyrt det kanvara att inte göra det. Att vara en skeptiker är att odla "street smarts" ikampen om kontrollen över sitt eget sinne, ens egna pengar, ett egetlojaliteter. För att vara en skeptiker, kort sagt, är att vägra att vara ett offer.- Robert S. DeBear "En agenda för Reason, realism och ansvar" New York Skeptic (nyhetsbrev New York området Skeptiker, Inc.), Spring 1988
		-- Cal Keegan

%
"Om du vill veta vad som händer med dig när du dör, gå titta på några dödagrejer."
		-- Dave Enyeart

%
"Efter en vecka [besöker Österrike] Jag kunde inte vänta med att gå tillbaka till FörentaStater. Allt var mycket trevligare i USA, på grund avmentalitet av att vara öppen, alltid positiv. Allt du villgöra i Europa är bara, "Inte en chans. Ingen har någonsin gjort det. " De har inte någonmer en önskan att gå ut för att erövra och uppnå - jag insåg att jag hade mycketmer den amerikanska andan. "
		-- Arnold Schwarzenegger

%
"Jag föredrar skurkar till idioter, eftersom de ibland ta en paus."
		-- Alexandre Dumas (fils)

%
Jag tror för det mesta att läsekretsen här använder c-ordet iett liknande sätt. Jag tror inte att någon verkligen tror på ett nytt, revolu-Ary litteratur --- Jag tror att de använder 'cyberpunk "som en term av bekvämlighetdiskutera gemensamma stilistiska element i en liten delmängd av de senaste sf böcker.
		-- Jeff G. Bone

%
Så vi får till min poäng. Visst folk häromkring läsa saker sominte på * officiellt sanktionerade Cyberpunk litteraturlista *. Visst viinte (någon av oss) verkligen tror att det finns några stora, djupa politiska ochfilosofiska budskap i allt detta, gör vi? Så om detta 'cyberpunk "sak ärbara en period av bekvämlighet, hur kan någon sälja ut? Om cyberpunk är bara enord vi använder för att beskriva en viss stil och bildspråk i sf, hur kan det varadöd? Var är den djupa uttalanden som det så kallade rörelsen "är eller försökteatt göra?Jag tror att de flesta av oss är intresserad av att undersöka och diskutera litterära(Och musikalisk) verk som besitter en viss stilistisk kvalitet och kanske enganska extrema perspektiv; detta är vad CP handlar om, eller hur? kanske finnsbör vara en diskussionsgrupp som, säg, alt.postmodern eller något. något mindrerestriktiv i omfattning än alt.cyberpunk.
		-- Jeff G. Bone

%
"Allas huvud är en billig film show."
		-- Jeff G. Bone

%
Livet är fullt av begrepp som är dåligt definierade. I själva verket finns det mycket fåbegrepp som inte är det. Det är svårt att tänka sig något i icke-tekniska områden.
		-- Daniel Kimberg

%
... Cyberpunk vill se sinnet som mekanistiska & duplicable,utmanande grundläggande antaganden om vilken typ av individualitet som själv.Det verkar allt bättre skäl att anta att cyberpunk konst & musik ärväsentligen mindless garbagio. Willy behandlas verkligen denna idé i"Count Zero" med Katatonenkunst den automatiska box-maker och flickansobservation att den verkliga konsten var byggandet av själva maskinen,snarare än dess utgång.
		-- Eliot Handelman

%
Det kan vara värt att reflektera att denna grupp skapades ursprungligentillbaka i september 1987 och har utväxlat över 1200 meddelanden. Deursprungliga meddelandet för grupp som kallas för en all inclusivediskussion som sträcker sig från handstilarna av Gibson och Vinge och filmersom Bladerunner till verkliga saker som Brands beskrivning avarbete som görs vid MIT Media Lab. Det var tänkt som en fristad förmänniskor med vision av denna omfattning. Om du vill skapa en fristad förpersoner med smalare visioner, gärna. Men jag känner mig ledsen för allasom tycker att alt.cyberpunk är en sådan monstruös grupp som det är iträngande behov av att delas. Heaven hjälpa dem om de någonsin startarläsning comp.arch eller rec.arts.sf-älskare.
		-- Bob Webber

%
... Jag bryr mig inte om begreppet "mekanistiska". Ordet "cybernetiska" är en mycketmer apropos. Den mekanistiska världsbilden faller allt längre bakomden verkliga världen där även enkla system kan producera de mest fantastiskakaos.
		-- Peter da Silva

%
När det gäller de grundläggande antaganden om individualitet och sig själv, är detta kärnanav vad jag tycker om cyberpunk. Och det är kärnan i vad jag tycker om vissapre-gibson neophile techie SF författare som vissa människor här vilja sättaner. Inte alla gör samma antaganden. Jag har inte förlorat mitt sinne ... det ärbackas upp på band.
		-- Peter da Silva

%
Vilka är konstnärerna i Computer Graphics Show? Wavefront senaste låda, ellerde människor som programmeras det? Skulle Mandelbrot få all kredit förproduktion av program som MandelVroom?
		-- Peter da Silva

%
Bakkant Technologies är glada att tillkännage följandeTETflame programmet:1) För en förhandlingslösning pris (inga quatloos accepteras) en av våra flammande   representanter flamma den levande skiten ur affischen av   ditt val. Priset är inversly proportionell mot hur mycket av   en skitstövel målet det. Vi kan inte vara övertygad om att flamma Dennis   Ritchie. Matt Crawford flammor är gratis.2) För en förhandlingslösning pris (samma arrangemang) den TETflame programmet   erbjuder `` flamma Insurence ''. Enligt detta arrangemang, om   en av våra försäkringstagare är flammade kommer vi avbryta den felande   artikeln och flamma den flamer, till en skarp.3) TETflame flammande representanter är: Richard Sexton, Oleg   Kisalev, Diane Holt, Trish O'Tauma, Dave Hill, Greg Nowak och vår mest   nyförvärv, Keith Doyle. Men allt han kommer att göra är att sätta dig i sitt   döda fil. Weemba enligt överenskommelse.
		-- Richard Sexton

%
"När jag gick bland bränder i Helvetet, glad med njutningar Geni; som till änglar ser ut som plåga och galenskap. Jag samlat några av deras Ordspråksboken ... "- Blake," Äktenskapet mellan himmel och helvete "
		-- Richard Sexton

%
HUR att bevisa det, DEL 1bevis med gott exempel:Författaren ger endast fallet n = 2 och antyder att detinnehåller de flesta av idéerna i den allmänna bevis.bevis genom hotelser:"Trivial".bevis genom kraftig handwaving:Fungerar bra i ett klassrum eller seminarium inställning.
		-- Richard Sexton

%
HUR att bevisa det, DEL 2bevis av besvärliga notation:Bäst med tillgång till minst fyra bokstäver och speciellasymboler.bevis genom utmattning:En fråga eller två av en tidskrift som ägnas åt ditt bevis är användbar.bevis genom utelämnande:"Läsaren kan lätt tillhandahålla detaljerna""De övriga 253 fall är analoga""..."
		-- Richard Sexton

%
HUR att bevisa det, DEL 3bevis av förvirring:En lång plotless sekvens av sann och / eller meningssyntaktiskt relaterade uttalanden.bevis av önske citat:Författaren citerar negationen, samtala, eller generalisering aven sats från litteraturen för att stödja sina påståenden.bevis av finansiering:Hur kunde tre olika myndigheter vara fel?bevis av framstående myndighet:"Jag såg Karp i hissen och han sade att det var förmodligen NPkomplett. '
		-- Richard Sexton

%
HUR att bevisa det, DEL 4bevis genom personlig kommunikation:"Åtta-dimensionell färgad cykel stripp är NP-komplett[Karp, personlig kommunikation]. "bevis genom reduktion till fel problem:"Att se att oändligt-dimensionell färgad cykel stripp äravgör minskar vi den till stopproblemet. "bevis med hänvisning till otillgängliga litteratur:Författaren citerar en enkel följd av en sats återfinnsi en privat cirkulerat memoar av den slovenskaFilologiska Society, 1883.bevis av betydelse:En stor mängd användbara konsekvenser alla följer avproposition i fråga.
		-- Richard Sexton

%
HUR att bevisa det, DEL 5bevis av ackumulerade bevis:Lång och omsorgsfull efterforskning har inte avslöjat en motexempel.bevis av kosmologin:Negationen av påståendet är otänkbart ellermeningslös. Populär för bevis för Guds existens.bevis genom ömsesidigt referens:Med hänvisning A, sats 5 sägs följa från Sats 3 ireferens B, som har visat sig följa från Korollarium 6,2 ireferens C, som är en enkel följd av Sats 5 ireferens A.bevis genom metaproof:En metod ges för att konstruera den önskade bevis. Dekorrekthet av metoden bevisas av någon av dessatekniker.
		-- Richard Sexton

%
HUR att bevisa det, DEL 6bevis för bild:En mer övertygande form av bevis med gott exempel. kombinerar bramed bevis genom utelämnande.yrkande genom häftig påstående:Det är bra att ha någon form av myndighet förhållande tillpublik.bevis genom spöke referens:Inget ens tillnärmelsevis liknar den citerade sats visas ireferensen.
		-- Richard Sexton

%
HUR att bevisa det, DEL 7bevis genom framåt referens:Referensen vanligtvis till ett kommande papper av författaren,vilket är ofta inte så kommande som i början.bevis av semantisk skift:Några av de vanliga men obekväma definitioner ändrasför redovisning av resultatet.bevis genom överklagande till intuition:Cloud-formade ritningar hjälpa ofta här.
		-- Richard Sexton

%
        [Maj en] tvivlar, i ost och trä, är maskar genereras,        eller, om skalbaggar och getingar, i ko-dynga, eller om fjärilar, gräshoppor,        skaldjur, sniglar, ål, och sådant liv att procreated av putrefied        materia, som skall motta formen av den varelsen till vilken den        är av formativ kraft anordnad [?] Att ifrågasätta detta är att ifrågasätta        Därför känsla och erfarenhet. Om han tvivlar detta, låt honom gå till        Egypten och där han hittar fält svärmar med möss födde        av leran av Nylus, till stor olycka av invånarna.                En sextonhundratalet yttrande citeras av L. L. Woodruff,                i * Utvecklingen av jorden och människan * 1929
		-- Richard Sexton

%
Sett på en knapp på en SF-konventionen:Veteran av Bermudatriangeln expeditionsstyrkan. 1990-1951.
		-- Richard Sexton

%
"Om människor är bra bara för att de är rädda för straff, och hoppas på belöning,då vi är en ledsen mycket faktiskt. "
		-- Albert Einstein

%
"Vad som önskas är inte viljan att tro, men viljan att ta reda på, vilket ärraka motsatsen. "
		-- Bertrand Russell, _Sceptical_Essays_, 1928

%
"Fanns det inga kvinnor, kan män leva som gudar."
		-- Thomas Dekker

%
"Intelligens utan tecken är en farlig sak."
		-- G. Steinem

%
"Det säger att han gjorde oss alla att vara precis som honom. Så om vi är dumma, är GUDstum, och kanske till och med lite ful på sidan. "
		-- Frank Zappa

%
"Det är inte bara en dator - det är din röv."
		-- Cal Keegan

%
"Låt mig gissa, Ed. Pentescostal, eller hur?"- Starcap'n Ra, ra@asuvax.asu.edu. "Nej karismatiska (jag tror - jag har gett upp vad alla de där irriterande etiketter betyda)."- Ed Carp, erc@unisec.usi.com"Samma skillnad - allt nit och känsla, i genomsnitt mindre än en arbetsdag hjärnacell per församling. Starcap'n Ra, knuten du honom. Bra jobbat!"
		-- Kenn Barry, barry@eos.UUCP

%
"BTW, inte Jesus vet du flamma?"
		-- Diane Holt, dianeh@binky.UUCP, to Ed Carp

%
"Jag har sett förfalskningar jag har skickats ut."
		-- John F. Haugh II (jfh@rpp386.Dallas.TX.US), about forging net news articles

%
"Bara av nyfikenhet betyder det faktiskt något eller har någon av de få återstående bitarna av din hjärna just avdunstat? "
		-- Patricia O Tuama, rissa@killer.DALLAS.TX.US

%
"Bite off, Dirtball."Richard Sexton, richard@gryphon.COM
		-- Patricia O Tuama, rissa@killer.DALLAS.TX.US

%
"Oh my! En` inflammatorisk attityd "i alt.flame? Aldrig hört talas om en sådanen sak..."
		-- Allen Gwinn, allen@sulaco.Sigma.COM

%
(Null kaka, hoppas det är ok)
		-- Allen Gwinn, allen@sulaco.Sigma.COM

%
"I kristendomen varken moral nor religion komma i kontakt med verklighetenvid någon punkt. "
		-- Friedrich Nietzsche

%
"Vem är ensam anledning att * ligga ut sig * av verkligheten? Han som * lider * från det."
		-- Friedrich Nietzsche

%
"Du som hatar judarna så, varför du anta sin religion?"
		-- Friedrich Nietzsche, addressing anti-semitic Christians

%
"Little prigs och trekvarts galningar kan ha inbilskhet att lagarna inatur ständigt bryts för deras skull. "
		-- Friedrich Nietzsche

%
"Vetenskapen gör godlike - det är hela med präster och gudar när man blir vetenskaplig. Moral: vetenskap är förbjuden som sådan - det enbart är förbjuden. Vetenskap är * första * synd, * ursprungliga * synd. * Bara detta är moral * `` Du skall inte vet '' -.. resten följer "
		-- Friedrich Nietzsche

%
"Tro: inte * vill * veta vad som är sant."
		-- Friedrich Nietzsche

%
> En grundläggande begrepp som ligger till grund Usenet är att det är ett kooperativ.Efter att ha varit på Usenet för att gå på tio år, jag håller inte med detta.Den grundläggande idén bakom Usenet är lågan.
		-- Chuq Von Rospach, chuq@Apple.COM

%
"Varje grupp har ett par experter. Och varje grupp har åtminstone en idiot. Således är balans och harmoni (och oenighet) upprätthålls. Det är ibland svårt att komma ihåg detta i huvuddelen av de e-gräl att alla besvär och smärta orsakas vanligtvis av en eller två högt motiverade, frätande twits. "
		-- Chuq Von Rospach, chuq@apple.com, about Usenet

%
Backas upp systemet på sistone?
		-- Chuq Von Rospach, chuq@apple.com, about Usenet

%
"Det är inte mycket beteckna som ett gifter för en är säker på att hitta ut nästamorgon det var någon annan. "
		-- Rogers

%
"Om du är rädd för ensamheten, inte gifta sig."
		-- Chekhov

%
"Love är en idealisk sak, äktenskapet en real thing, en sammanblandning av den verkliga medden ideala går aldrig ostraffad. "
		-- Goethe

%
"I äktenskap, att tveka ibland ska sparas."
		-- Butler

%
"Den stora frågan ... som jag inte har kunnat svara ... är, 'Vad görkvinna vill ha? ""
		-- Sigmund Freud

%
"Jag har nyligen undersökt alla de kända vidskepelserna av världen, och inte hittar i vår särskilda vidskepelse (kristendomen) en försonande särdrag. De är alla lika bygger på fabler och mytologi. "
		-- Thomas Jefferson

%
Kom ihåg: Silly är ett sinnestillstånd, är dumma ett sätt att leva.
		-- Dave Butler

%
"The främste av en lärd man över en dyrkare är lika med den främsteav månen, på natten av fullmånen, över alla stjärnor. Sannerligen, denlärda män är arvtagare av profeterna. "
		-- A tradition attributed to Muhammad

%
"The präster framgångsrikt predikade läror tålamod och pusillanimity;de aktiva dygderna i samhället har avskräckt; och de sista resterna av enmilitär anda begravdes i klostret: en stor del av allmänheten ochprivat rikedom invigdes till bestickande krav välgörenhet och hängivenhet;och soldaternas löner var får på onödiga mängder av båda könensom bara kunde åberopa fördelarna med avhållsamhet och kyskhet. "
		-- Edward Gibbons, _The Decline and Fall of the Roman Empire_

%
"Frågan är snarare: om vi någonsin lyckas göra ett sinne" nötterbultar ", hur ska vi vet att vi har lyckats?- Fergal Toomey"Det kommer att berätta."
		-- Barry Kort

%
"Förfrågan är dödlig till visshet."
		-- Will Durant

%
"Mets var stor i" sextioåtta, Korten var bra i "sextio nio, Men lejonungarna kommer att bli himmelsk i nitton och sjuttio. "
		-- Ernie Banks

%
"Vid två tillfällen jag har blivit ombedd [av riksdagsledamöter!]," Be, Mr.Babbage, om du sätter in i maskinen fel siffror, kommer de rätta svarenkomma ut?' Jag kan inte riktigt att uppfatta den typ av begreppsförvirringsom kan framkalla en sådan fråga. "
		-- Charles Babbage

%
"Jag kallar kristendomen * en * stor förbannelse, det * en * stor inneboendefördärv, det * en * bra instinkt för hämnd för vilken ingen utvägär tillräckligt giftig, hemlig, underjordisk, * småaktiga * - Jag kallar det* Ett * dödlig fläck för mänskligheten. "
		-- Friedrich Nietzsche

%
"Det grundläggande syftet animera Guds Tro och Hans religion är atttillvarata och främja enighet av mänskligheten, och för att främjaen anda av kärlek och gemenskap bland män. Lider det inte att bli en källaav oenighet och oenighet, hat och fiendskap. ""Religionen är sannerligen huvudinstrumentet för att inrätta ordning i värld och lugn bland det folk ... Ju större nedgång religion, desto mer smärtsamma den egensinnighet av de ogudaktiga. Detta kan inte annat än bly i slutet för att kaos och förvirring. "
		-- Baha'u'llah, a selection from the Baha'i scripture

%
"Cogito ergo jag har rätt och du har fel."
		-- Blair Houghton

%
"... En av de främsta orsakerna till nedgången av det romerska riket var attsaknar noll, hade de inget sätt att indikera framgångsrik avslutning avderas C-program. "
		-- Robert Firth

%
Q: Någon precis postat att Roman Polanski riktade Star Wars. Vadborde jag?A: Skicka rätt svar på en gång! Vi kan inte ha folk gå på troden där! Mycket bra av dig att upptäcka detta. Du kommer förmodligen att vara den enda somgöra korrigeringen, så skicka så fort som möjligt. Ingen tid att förlora, såverkligen inte vänta en dag, eller kontrollera om någon annan har gjortkorrektion.Och det är inte tillräckligt bra för att skicka meddelandet per post. Eftersom du är denenda som verkligen vet att det var Francis Coppola, du måste informerahela nätet direkt!
		-- Brad Templeton, _Emily Postnews Answers Your Questions on Netiquette_

%
Fråga: Hur kan jag välja vilka grupper för att skriva in? ...Fråga: Hur ett exempel?A, okej. Låt oss säga att du vill rapportera att Gretzky har handlats frånOilers till Kings. Nu genast du kanske tror rec.sport.hockeyskulle vara tillräckligt. FEL. Många fler människor kan vara intresserade. Det här är enstor handel! Eftersom det är en nyhetsartikel, hör det i nyheterna. * Hierarkinockså. Om du är en nyhets admin, eller om det finns en på din dator, försöknews.admin. Om inte, använd news.misc.De Oilers är förmodligen intresserad av geologi, så försök sci.physics. Han ären stor stjärna, så skicka till sci.astro och sci.space eftersom de är ocksåintresserad av stjärnor. Därefter är hans namn polska klingande. Så skicka tillsoc.culture.polish. Men den gruppen inte existerar, så kors post tillnews.groups tyder det bör skapas. Med så här många grupper avintresse, kommer din artikel vara ganska bisarra, så skicka till talk.bizarre somväl. (Och lägga till comp.std.mumps, eftersom de knappast få några artiklardär, och en "comp" grupp kommer att fortplanta din artikel ytterligare.)Du kan också finna det är roligare att skriva artikeln en gång i varje grupp.Om du lista alla diskussionsgrupper i samma artikel, några diskussionsgruppsläsare kommerendast visar artikeln för att läsaren en gång! Inte tolerera detta.
		-- Brad Templeton, _Emily Postnews Answers Your Questions on Netiquette_

%
Fråga: Jag kan inte stava värd en fördämning. Jag hoppas du kommer också säga vad jag ska göra?A: Bry dig inte om hur dina artiklar ser ut. Kom ihåg att det är meddelandetsom räknas, inte hur det presenteras. Bortse från det faktum att slarvigastavningen i ett helt skriftligt forum sänder ut samma tysta meddelanden somnedsmutsade kläder skulle när man behandlar en publik.
		-- Brad Templeton, _Emily Postnews Answers Your Questions on Netiquette_

%
Q: De meddelade bara på radion att Dan Quayle valdes somRepublikan V.P. kandidat. Ska jag lägga?A: Självklart. Nätet kan nå människor på så lite som 3-5 dagar. Dessdet perfekta sättet att informera om sådana nyhetshändelser långt efterbroadcast nätverk har täckt dem. Som ni förmodligen den enda personenatt ha hört nyheten på radion, vara noga med att lägga så fort som möjligt.
		-- Brad Templeton, _Emily Postnews Answers Your Questions on Netiquette_

%
Vad gjorde Mickey Mouse få till jul?En Dan Quayle klocka.
		-- heard from a Mike Dukakis field worker

%
Fråga: Vad är skillnaden mellan en bilförsäljare och en dator    försäljare?A: bilförsäljare kan förmodligen köra!
		-- Joan McGalliard (jem@latcs1.oz.au)

%
"Din dumhet, Allen, är helt enkelt inte upp till par."- Dave Mack (mack@inco.UUCP)"Yours är."
		-- Allen Gwinn (allen@sulaco.sigma.com), in alt.flame

%
Ett urval av de taoistiska skrifter:"Lao-Tan frågade Konfucius: 'Vad menar du med välvilja och rättfärdighet"? Konfucius sade: 'Att vara i sitt innersta hjärta i vänligt sympati med alla saker; att älska alla män och låta några själviska tankar: det är naturen av välvilja och rättfärdighet. ' "
		-- Kwang-tzu

%
"Jesus sparar ... men Gretzky får rebound!"
		-- Daniel Hinojosa (hinojosa@hp-sdd)

%
"Allt som skapats måste med nödvändighet vara sämre än kärnan i skaparen."- Claude Shouse (shouse@macomw.ARPA)"Einsteins mamma måste ha varit ett fan av en fysiker."
		-- Joseph C. Wang (joe@athena.mit.edu)

%
"Religionen är något kvar från barndom vår intelligens, det kommerblekna bort som vi antar skäl och vetenskap som våra riktlinjer. "
		-- Bertrand Russell

%
"Lögnaktiga läppar är en styggelse för Herren, men de som handlar verkligen är hans glädje. Ett mjukt svar stillar vrede; men ord som sårar väcker ilska. Han som svarade en fråga innan han hör det, är det dårskap och skam till Hej M. Inte vara en vittnesbörd mot din nästa utan sak; och lura inte med dina läppar. Död och liv är i kraft av tungan. "
		-- Proverbs, some selections from the Jewish Scripture

%
"Som en tonåring jag strävat efter att varaktig berömmelse, längtade jag faktisk säkerhet, ochJag törstade efter en meningsfull vision av mänskligt liv - så jag blev en vetenskapsman.Detta är som att bli en ärkebiskop så att du kan träffa tjejer. "
		-- Matt Cartmill

%
Heisenberg kan ha varit här.
		-- Matt Cartmill

%
"Någon ursäkt kommer att tjäna en tyrann."
		-- Aesop

%
"Erfarenheten har visat att vissa människor verkligen vet allt."
		-- Russell Baker

%
Hur många Zenbuddist tar det att byta en glödlampa?Två. En ändra det och en inte att ändra det.
		-- Russell Baker

%
"Jag föredrar trubbiga påkar av anhängarna av ormen Gud."
		-- Sean Doran the Younger

%
"Om jag inte vill att andra ska citera mig, jag talar inte."
		-- Phil Wayne

%
"Min terminal är en dödlig tesked."
		-- Patricia O Tuama

%
"Jag är ... en kvinna ... och ... tekniskt en parasitisk livmodertillväxt"
		-- Sean Doran the Younger [allegedly]

%
"Är det bara jag, eller är det någon annan läsa` bibel Humpers "varje gångnågon skriver 'bibel thumpers?
		-- Joel M. Snyder, jms@mis.arizona.edu

%
"Pengar är roten till allt pengar."
		-- the moving finger

%
"... Greg Nowak: 'En annan lågan från Greg" - behöver jag säga mer? "- Jonathan D. Trudel, trudel@caip.rutgers.edu"Nej, du måste säga mindre."
		-- Richard Sexton, richard@gryphon.COM

%
"Och det är min åsikt, och det är bara min åsikt, du är en galning. Justeftersom det inte finns några hunderd andra personer som delar din vansinne med diggör dig inte någon sundare. Dömd, va? "
		-- Oleg Kiselev,oleg@CS.UCLA.EDU

%
"Lydnad. En religion av slavar. En religion av intellektuell död. Jag gillarDet. Inte ställa frågor, tror inte, lyder Herrens ord - som dethar bekvämt lett till dig av en man i en Rolls med en tung Rolexpå hans handled. Jag gillar det jobbet! Var kan jag registrera? "
		-- Oleg Kiselev,oleg@CS.UCLA.EDU

%
"Home liv som vi förstår det är inte mer naturligt för oss än en bur är att enkakadua."
		-- George Bernard Shaw

%
"Äktenskapet är som en bur, man ser fåglarna utanför desperat att komma in, ochde inne desperata att komma ut. "
		-- Montaigne

%
"För en manlig och kvinnlig leva kontinuerligt tillsammans är ... biologisktsett en extremt onaturligt tillstånd. "
		-- Robert Briffault

%
"Äktenskapet är lågt, men du tillbringa resten av ditt liv att betala för det."
		-- Baskins

%
En man är inte komplett förrän han är gift - då han är klar.
		-- Baskins

%
Äktenskapet är den enda orsaken till skilsmässa.
		-- Baskins

%
Äktenskapet är en triumf för fantasin över intelligens. Andra äktenskap ärden hoppets triumf över erfarenheten.
		-- Baskins

%
"Kedjan som kan slet är inte den eviga kedjan."
		-- G. Fitch

%
"Gå till himmel för klimatet, helvete för företaget."
		-- Mark Twain

%
"Jag är övertygad om att tillverkarna av matt ta bort lukt pulver har ingår inkapslade tid släpptes katt urin i sina produkter. Detta teknik måste vara vad hindrade dess fördelning under min mammas regeringstid. Min Mattan luktar piss och jag har inte en katt. Bättre gå med lite mer. "
		-- timw@zeb.USWest.COM, in alt.conspiracy

%
"Om det inte finns en befolkning problem, varför är regeringen att sätta cancer icigaretterna? "
		-- the elder Steptoe, c. 1970

%
"Om du inte vill att din hund att ha dålig andedräkt, gör vad jag: Häll lite Lavoris i toaletten. "
		-- Comedian Jay Leno

%
"Här är något att tänka på: Hur kommer du aldrig se en rubrik som `Psychic vinner lotteri."
		-- Comedian Jay Leno

%
"Well hello there Charlie Brown, fåntratt dig."
		-- Lucy Van Pelt

%
"Time är en illusion. Lunchtid dubbelt så."
		-- Ford Prefect, _Hitchhiker's Guide to the Galaxy_

%
"Okunnighet är jorden där tron ​​på mirakel växer."
		-- Robert G. Ingersoll

%
"Låt var och en lära sin son, lära sin dotter, att arbetet är hedervärd."
		-- Robert G. Ingersoll

%
"Jag har inte den minsta tilltro till" andliga manifestationer. "
		-- Robert G. Ingersoll

%
"Det är svårt att överskatta den skuld som vi är skyldiga att män och kvinnor i geni."
		-- Robert G. Ingersoll

%
"Joy är rikedom och kärlek är lagligt betalningsmedel i själen."
		-- Robert G. Ingersoll

%
"Händerna som hjälper är bättre långt än läpparna som ber."
		-- Robert G. Ingersoll

%
"Det är kreationist som hädiskt hävdar att Gud fusk oss på ett dumt sätt. "
		-- J. W. Nienhuys

%
"Nej, nej, jag inte emot att kallas den smartaste mannen i världen. Jag önskar bara det inte var här. "
		-- Adrian Veidt/Ozymandias, WATCHMEN

%
"Var * utmärkt * till varandra."
		-- Bill, or Ted, in Bill and Ted's Excellent Adventure

%
Den sjunde upplagan tillståndsförfaranden är, antar jag, fortfarande i kraft,även om jag tvivlar på att band är tillgängliga från AT & T. I varje fall, oberoenderestriktioner licensen ställer fortfarande existerar. Dessa begränsningar var ochär rimliga för platser som bara vill köra systemet, men tillåter intemånga av de saker som Minix skrevs för, liksom studier av källan iklasser, eller av personer som inte på ett universitet eller företag.Jag har alltid trott att Minix var en fin idé, och kompetent gjort.Som för storleken på v7, wc -l /usr/sys/*/*.[chs] är 19.271.
		-- Dennis Ritchie, 1989

%
"Vår vision är att påskynda tid, så småningom eliminera det." - Alex Schure
		-- Dennis Ritchie, 1989

%
"Kärlek är en snöskoter racing över tundra och sedan plötsligt flippar över, sätter du nedanför. På natten, isen vesslor komma. "
		-- Matt Groening

%
"Jag är inte rädd för att dö, jag vill bara inte att vara där när det händer."
		-- Woody Allen

%
"The Street finner sina egna användningsområden för tekniken."
		-- William Gibson

%
"Jag ser lite gudomlighet om dem eller dig. Du pratar med mig om kristendomennär du är i färd med att hänga dina fiender. Fanns det någonsin en sådanhädiska nonsens! "
		-- Shaw, "The Devil's Disciple"

%
"Du och jag som individer kan genom upplåning, leva över våra tillgångar, menbara under en begränsad tid. Varför ska vi tro att kollektivt,som en nation, vi är inte bundna av samma begränsning? "
		-- Ronald Reagan

%
"Han gjorde besluta om att med mer tid och en hel del mental ansträngning,han skulle förmodligen vända verksamheten till en acceptabel perversion. "
		-- Mick Farren, _When Gravity Fails_

%
"Konvertering, sparsmakad gudinna, älskar blod bättre än tegel och festermest subtilt på den mänskliga viljan. "
		-- Virginia Woolf, "Mrs. Dalloway"

%
Det är dags att starta upp, gör din boot rom vet var dina diskkontroller är?
		-- Virginia Woolf, "Mrs. Dalloway"

%
"Vad forskarna har i sina portföljer är skrämmande."
		-- Nikita Khrushchev

%
"... En mest utmärkta barbar ... Djingis Kahn!"
		-- _Bill And Ted's Excellent Adventure_

%
"Tryck på avtryckaren och du är skräp."
		-- Lady Blue

%
"Åh vad skulle jag inte ge vara spottade på i ansiktet ..."
		-- a prisoner in "Life of Brian"

%
"Sanningen aldrig kommer till världen men som en oäkting, till smälekav honom som förde hennes födelse. "
		-- Milton

%
"Om du inte kan debattera mig, då finns det inget sätt i helvetet du out-förolämpa mig."- Scott Legrand (Scott.Legrand@hogbbs.Fidonet.Org)"Du kan ha fel här, lilla."
		-- R. W. F. Clark (RWC102@PSUVM)

%
"Ja, jag är en verkligt arbete. En sak som vi lär sig ULowell är hur man flamma värdelös dataintrång icke-EE är som du. Jag är överlägsen dig i alla sätt genom utbildning och kompetens inom det tekniska området. Vem som helst kan lära sig hur man hacka, men teknik kommer inte alls lika lätt. Egentligen är jag inte försöker förolämpa alla du CS majors där ute, men jag tror EE är en av de svåraste majors / grad stora företagen att passera. Lyckligtvis, jag gör det. "- "Warrior Diagnostics" (wardiag@sky.COM)"Att både en EE och en skitstövel samtidigt måste vara en fruktansvärd börda till dig. Detta är egentligen inte en flamma, bara en tillfällig observation. Gör mig glad att jag var en CS major, livet är riktigt trevlig för mig. Ha kul med din valda läget av existens! "
		-- Jim Morrison (morrisj@mist.cs.orst.edu)

%
"BYTE redaktörer är män som skiljer agnarna från vetet, och sedan ut vetet. "
		-- Lionel Hummel (uiucdcs!hummel), derived from a quote by Adlai Stevenson, Sr.

%
DEN "FUN WITH USENET" MANIFESTMycket lite händer på Usenet utan någon form av svar från någon annanläsare. Fun With Usenet inlägg är inget undantag. Eftersom det finns några somkan ifrågasätta den logiska grunden för vissa av de utdrag som ingår däri, har jagskrivs en lista med riktlinjer som sammanfattar filosofin bakom dessainlägg.	En. Jag skar aldrig ut ord i mitten av ett citat utan en mycketgoda skäl, och jag skär dem aldrig utan inklusive ellipser. Förexempel: "Jag är inte en goob" kan bli "Jag är ... en goob", men det är ocksåvardagliga bry sig. "Jag är flamsäker" kan (och har) blir"Jag är ... en ... p ... oof", men det är verkligen sträcker sig det.Två. Om jag skär ord utanför början eller slutet av en offert, gör jag intesätta ellipser, men inte heller jag kapitalisera något som inte var aktiveradeinnan snittet. "Jag tror inte att kyrkan Ubizmo är en underbarplats "skulle förvandlas till" kyrkan Ubizmo är en underbar plats ". Tänkutstationering som en bandinspelning av affischen tankar. Om jag kan ställaupp citatet via snabbspola framåt och stoppa bandet, och utan splitsning,Jag lägger inte ellipser i. Och förresten, jag älskar att använda denna mekanism förvrida saker runt. Om du tror att något stinker, säger så - säg inte att dutror inte att det är underbart. ...
		-- D. J. McCarthy (dmccart@cadape.UUCP)

%
"De som kan ge upp nödvändig frihet att erhålla en lite tillfälligsäkerhet förtjänar varken frihet eller säkerhet. "
		-- Benjamin Franklin, 1759

%
"Jag är därför jag är."
		-- Akira

%
"Stan och jag trodde att detta experiment var så dum, beslutade vi att finansiera det själva. "
		-- Martin Fleischmann, co-discoverer of room-temperature fusion (?)

%
"Jag har mer information på ett ställe än någon i världen."
		-- Jerry Pournelle, an absurd notion, apparently about the BIX BBS

%
"Det är vad du lär när du vet allt som räknas."
		-- John Wooden

%
#define BITCOUNT (x) (((BX_ (x) + (BX_ (x) >> 4)) & 0x0F0F0F0F)% 255)#define BX_ (x) ((x) - (((x) >> 1) & 0x77777777) \- (((X) >> 2) & 0x33333333) \- (((X) >> 3) & 0x11111111))
		-- really weird C code to count the number of bits in a word

%
"Om du kan skriva en nations berättelser, behöver du inte oroa dig som gör sin lagar. Idag, berättar tv flesta historier att de flesta människor större delen av tiden. "
		-- George Gerbner

%
"Den rimliga man anpassar sig till världen, den orimliga en kvarstår för att försöka anpassa världen med sig själv. Därför måste alla framsteg beror på orimligt mannen. "
		-- George Bernard Shaw

%
"Vi vill skapa dockor som drar sina egna strängar."- Ann Marion"Skulle detta gör dem marionett?"
		-- Jeff Daiell

%
När det gäller C-program indrag:"I min Egotistical yttrande, bör de flesta människors C-program vara indragen sex fot nedåt och täckt med smuts. "
		-- Blair P. Houghton

%
Det fanns, det dök upp, en mystisk rit om inledande genom vilken, iett eller annat sätt, nästan varje medlem i teamet passerat. Den term somde gamla händer som används för denna rit - West uppfann sikt inte praxis -var `registrerar dig." Genom att registrera dig för projektet som du gick med på att göra vad som helstvar nödvändigt för framgång. Du gick med på att överge, om så är nödvändigt, familj,hobbies, och vänner - om du haft något av dessa kvar (och du kanske inte, omdu hade skrivit upp för många gånger tidigare).
		-- Tracy Kidder, _The Soul of a New Machine_

%
"När de hade minskat från 50 till 8, började de andra dvärgarnaatt misstänka "Hungry".
		-- a Larson cartoon

%
"Men tror du inte kan färgen på vin i ett kristallglas vara andlig. Utseendet på ett ansikte, musik av en fiol. A Paris teater kan ges med det andliga för all sin soliditet. "
		-- Lestat, _The Vampire Lestat_, Anne Rice

%
"Älska ditt land, men aldrig lita på sin regering."
		-- from a hand-painted road sign in central Pennsylvania

%
      Jag köpte den senaste dator;      det kom fullastad.      Det garanteras för 90 dagar,      men i 30 var omoderna!
		-- The Wall Street Journal passed along by Big Red Computer's SCARLETT

%
För att uppdatera Voltaire: "Jag kan döda alla medd från dig, men jag ska kämpa fördin rätt att lägga upp den, och jag ska låta det ligga på mina diskar ".
		-- Doug Thompson (doug@isishq.FIDONET.ORG)

%
"Även om ett program, men tre rader lång,dag det kommer att finnas kvar. "
		-- The Tao of Programming

%
"Turn on, tune upp, rocka loss."
		-- Billy Gibbons

%
         JORD     smog | tegelstenar AIR - lera - FIREsodavatten | tequila         VATTEN
		-- Billy Gibbons

%
"Naturligtvis elverktyg och alkohol hör inte ihop. Alla vet elverktyg är intelösliga i alkohol ... "
		-- Crazy Nigel

%
"Livet suger, men döden inte släcka alls ...."
		-- Thomas J. Kopp

%
   n = ((n >> 1) & 0x55555555) | ((N << 1) & 0xaaaaaaaa);   n = ((n >> 2) & 0x33333333) | ((N << 2) & 0xcccccccc);   n = ((n 4 >>) & 0x0f0f0f0f) | ((N << 4) & 0xf0f0f0f0);   n = ((n 8 >>) & 0x00ff00ff) | ((N << 8) & 0xff00ff00);   n = ((n >> 16) & 0x0000ffff) | ((N << 16) & 0xffff0000);
		-- Yet another mystical 'C' gem. This one reverses the bits in a word.

%
"Överallt, från populärkulturen till propagandan systemet finns detkonstant tryck för att få folk att känna att de är hjälplösa, att den enda rollde kan ha är att ratificera beslut och att konsumera. "
		-- Noam Chomsky

%
"Ett komplext system som fungerar är alltid visade sig ha utvecklats från en enkelsystem som fungerade. "
		-- John Gall, _Systemantics_

%
"Enligt min mening, Richard Stallman skulle inte känna igen terrorism om detkom upp och bet honom på hans Internet. "
		-- Ross M. Greenberg

%
Jag gjorde det till en regel att underlåta alla direkta motsägelser till känslor avandra, och alla positiva påstående om min egen. Jag förbjöd även själv användningenvarje ord eller uttryck i språk som importerat en fast åsikt,såsom "säkert", "utan tvekan", etc. Jag antog i stället för dem "Itänka "," Jag uppfattar ", eller" Jag kan tänka mig "en sak att vara så eller så, eller" så detförefaller för närvarande ".När en annan hävdade något som jag trodde fel, förnekade jag självnöjet att motsäga honom plötsligt, och att visa honom omedelbart någraabsurditet i hans förslag. För att besvara började jag med att konstatera att ivissa fall eller omständigheter hans åsikt skulle vara rätt, men i dettafall föreföll eller tycktes mig en viss skillnad, etc.Jag fann snart fördelen med denna förändring i mitt sätt; samtalen Ibedriver gick på mer positivt. Den blygsamma sätt som jag föreslog minyttranden skaffade dem en mer redo mottagning och mindre motsägelse. jag hademindre förtret när jag befanns vara i fel, och jag lättaresegrade med andra för att ge upp sina misstag och gå med mig när jagråkade vara på rätt.
		-- Autobiography of Benjamin Franklin

%
"Om jag någonsin komma runt att skriva detta språk depompisifier, kommer det att förändranästan alla förekomster av ordet "paradigm" i "exempel" eller "modell".
		-- Herbie Blashtfalt

%
"Livet, avsky den eller ignorera det, du kan inte ha det."
		-- Marvin the paranoid android

%
Förakt ljus blixtrade över datorns konsol.
		-- Hitchhiker's Guide to the Galaxy

%
"Det måste vara ett misstag", sade han, "är du inte en större dator änden miljarder svenska Gargantubrain som kan räkna alla atomer i en stjärna i enmillisekund? ""The miljarder svenska Gargantubrain?" sade Deep Thought med ohöljd förakt."Enbart kulram. Nämn det inte."
		-- Hitchhiker's Guide to the Galaxy

%
"Men är du inte", sade han, "en mer djävulsk tvist än den stora HyperlobicOmni-besläktad Neutron Wrangler av Ciceronicus Tolv, Magic ochOuttröttlig?""The Great Hyperlobic Omni-besläktade Neutron Wrangler", säger djupa tankar,noggrant rulla R, "kunde tala alla fyra benen av en ArcturanMega-Donkey - men bara jag kunde förmå det att gå en promenad efteråt ".
		-- Hitchhiker's Guide to the Galaxy

%
Om byggare byggde byggnader vägen programmerare skriver program, Jolt Colaskulle vara ett Fortune-500 företag.Om byggare byggde byggnader vägen programmerare skriver program, skulle du varakunna köpa en fin liten koloniala etage på Babbages för $ 34,95.Om programmerare skrev program vägen byggare bygga hus, skulle vi fortfarandevara att använda autocoder igång Samla däck.
		-- Peter da Silva and Karl Lehenbauer, a different perspective

%
Att fela är mänskligt, att moo nötkreatur.
		-- Peter da Silva and Karl Lehenbauer, a different perspective

%
"Amerika är en starkare nation för ACLU kompromisslösa ansträngning."
		-- President John F. Kennedy

%
"De enkla rättigheter, medborgerliga friheter från generationer av kamp får intebli bra ord för patriotiska semester, ord som vi undergräva på vardagar, menlevande, hedrade uppföranderegler bland oss ​​... Jag är glad att det amerikanska inbördesLiberties Union blir indignerad, och jag hoppas att detta kommer alltid att vara så. "
		-- Senator Adlai E. Stevenson

%
"Den ACLU har stått fyrkant mot de återkommande tidvatten av hysteri somfrån tid till annan hotar friheter överallt ... I själva verket är det svårtatt uppskatta hur långt våra friheter kan ha eroderat det inte hade varit för denEU: s tapper representation vid domstol i de konstitutionella rättighetermänniskor av alla övertygelser, oavsett hur impopulär eller ens föraktadeav majoriteten de var vid den tiden. "
		-- former Supreme Court Chief Justice Earl Warren

%
"Styrkan i konstitutionen ligger helt i fastställandet av varjemedborgare för att försvara det. Endast om varje enskild medborgare känner skyldig att görasin andel i detta försvar är konstitutionella rättigheter säkra. "
		-- Albert Einstein

%
"Jo jag förstår inte varför jag måste göra en man olycklig när jag kan göra så mångamän lycklig. "
		-- Ellyn Mustard, about marriage

%
"Och det borde vara lag: Om du använder ordet 'paradigm" utan att veta vadordlistan säger att det betyder, du går till fängelse. Inga undantag."
		-- David Jones @ Megatest Corporation

%
"Luke, jag är yer pappa, va. Kom över till den mörka sidan, hoser dig."
		-- Dave Thomas, "Strange Brew"

%
"Låt oss inte vara alltför hårda på vår egen okunnighet. Det är det som gör Amerika stor. Om Amerika inte var ojämförligt okunniga, hur kunde vi har tolererat de senaste åtta åren? "
		-- Frank Zappa, Feb 1, 1989

%
"Historien om alla större Galactic Civilization tenderar att passera igenomtre distinkta och igenkännbara faser, de Överlevnad, Förfrågan ochFörfining, annars känd som hur, varför och var faser."Till exempel är den första fasen kännetecknas av frågan" Hur kanvi äter?' den andra av frågan "Varför äter vi?" och den tredje avfrågan "Var ska vi äta lunch?"
		-- Hitchhiker's Guide to the Galaxy

%
"Tro inte, låt maskinen göra det åt dig!"
		-- E. C. Berkeley

%
"Härav följer att någon överbefälhavare som åtar sig att genomföra en plan som han anser defekt är fel; han måste lägga fram sina skäl, insistera av planen ändras, och slutligen entledigande snarareän vara instrumentet för hans armé undergång. "
		-- Napoleon, "Military Maxims and Thought"

%
"(Chief programmerare) personligen definierar den funktionella och prestanda specifikationer, designar programmet, koder det, testar den, och skriver sin dokumentation ... Han behöver stor talang, tio års erfarenhet och avsevärda system och applikationer kunskap, vare sig i tillämpad matematik, affärsdata hantering, eller vad som helst. "
		-- Fred P. Brooks, _The Mythical Man Month_

%
"Det är inte över förrän det är över."
		-- Casey Stengel

%
"Om något kan gå fel, kommer det."
		-- Edsel Murphy

%
"Yo barn yo barn yo."
		-- Eddie Murphy

%
"Du måste lära dig att köra din kajak genom ett slags ju-jitsu. Du måste lära dig att berätta vad floden kommer att göra för dig, och med tanke på dessa parametrar se hur du kan leva med det. Du måste absorbera sin kraft och omvandla den till användarna så gott du kan. Även med snabbhet och smidighet i en kajak, du är inte snabbare än floden, eller starkare, och du kan slå det endast genom förstå den. "
		-- Strung, Curtis and Perry, _Whitewater_

%
Alla som kommer in här vill tre saker:1. De vill det snabbt.2. De vill ha det bra.3. De vill ha det billigt.Jag berättar dem att plocka två och ringa mig tillbaka.
		-- sign on the back wall of a small printing company in Delaware

%
"Fler mjukvaruprojekt har gått snett på grund av kalendertiden än för alla andra orsaker kombineras. "
		-- Fred Brooks, Jr., _The Mythical Man Month_

%
panik: kernel trap (ignoreras)
		-- Fred Brooks, Jr., _The Mythical Man Month_

%
"Kärnvapenkrig kan förstöra hela din kompilering."
		-- Karl Lehenbauer

%
"Kom ihåg, extremism i nondefense av moderation är inte en dygd."
		-- Peter Neumann, about usenet

%
"Vi ägnat oss till en kraftfull idé - organisk lag snarare än naken driva. Det verkar vara universell acceptans av denna idé i nationen. "
		-- Supreme Court Justice Potter Steart

%
"Vad man har gjort, kan man strävar efter att göra."
		-- Jerry Pournelle, about space flight

%
"Om du kan, hjälpa andra. Om du kan inte, åtminstone inte skadar andra."
		-- the Dalai Lama

%
Till system programmerare, användare och applikationer tjänar bara för att ge enprovbelastningen.
		-- the Dalai Lama

%
"Tänk, med VLSI vi kan ha 100 ENIACS på ett chip!"
		-- Alan Perlis

%
"... Lokala förbud kan inte blockera framsteg inom militära och kommersiella teknik ... demokratiska rörelser för lokal återhållsamhet kan bara hålla världens demokratier, inte världen som helhet. "
		-- K. Eric Drexler

%
"Den rotter som simpers att han ser ingen skillnad mellan en fem-dollarsedeloch en piska förtjänar att lära sig skillnaden på sin egen rygg - som, tror jag, hankommer."
		-- Francisco d'Anconia, in Ayn Rand's _Atlas Shrugged_

%
"Om en nation värderar något mer än frihet, kommer den att förlora sin frihet, och ironin av det är att om det är komfort eller pengar det värderar mer, kommer det förlora det också. "
		-- W. Somerset Maugham

%
"Förlåt mig för att andas, som jag aldrig göra hur som helst så jag vet inte varför jag bry att säga det, o Gud, jag är så deprimerad. Här är en annan av de självbelåten dörrar. Liv! Inte prata med mig om livet. "
		-- Marvin the Paranoid Android

%
En av de största svårigheterna Trillian upplevt i hennes relation medZaphod lärde sig att skilja mellan honom låtsas vara dum baraatt få människor utanför sin vakt, låtsas vara dum eftersom han inte kundevara störd att tänka och ville ha någon annan att göra det för honom, låtsasatt vara så skandalöst dumt att dölja det faktum att han faktiskt inte förståhatt pågick, och verkligen är genuint dum. Han var renowned förär ganska smart och helt klart var så - men inte hela tiden, vilketuppenbarligen oroade honom, därav lagen. Han föredrog folk att vara förbrylladsnarare än förakt. Detta framför allt tycktes Trillian att varagenuint dum, men hon kunde inte längre vara störd att argumentera om.
		-- Douglas Adams, _The Hitchhiker's Guide to the Galaxy_

%
Långt tillbaka i dimma gamla tiden, i de stora och härliga dagar itidigare Galactic Empire, var liv vild, rik och till stor del skattefria.Mäktiga rymdskepp levererat sin väg mellan exotiska solar, söker äventyr ochbelöna bland de längst når i Galactic utrymme. I dessa dagar, spritvar modig, insatserna var höga, män var riktiga män, kvinnor var riktiga kvinnoroch små lurviga varelser från Alpha Centauri var verkliga små lurviga varelserfrån Alpha Centauri. Och alla vågade trotsa okända skräck, att göra mäktiggärningar, att frimodigt dela infinitiv att ingen människa hade spruckit tidigare - och därmedvar Empire förfalskade.
		-- Douglas Adams, _The Hitchhiker's Guide to the Galaxy_

%
"Gort, Klaatu Nikto Barada."
		-- The Day the Earth Stood Still

%
> Från MAILER-DAEMON@Think.COM Thu 2 mars 13:59:11 1989> Ämne: Åter post: okänt mailer error 255"Dale, din adress inte längre fungerar. Kan du fixa det på din sida?"- Bill Wolfe (wtwolfe@hubcap.clemson.edu)"Bill, hjärnan inte längre fungerar. Kan du fixa det på din sida?"
		-- Karl A. Nyberg (nyberg@ajpo.sei.cmu.edu)

%
"Tappa inte syra, ta det pass-misslyckas!"
		-- Bryan Michael Wendt

%
"Jag fick en fråga för dig. Ya fick en minut?"
		-- two programmers passing in the hall

%
Jag tog en fisk huvud på bio och jag behövde inte betala.
		-- Fish Heads, Saturday Night Live, 1977.

%
Vad har Bob åstadkommit?
		-- Fish Heads, Saturday Night Live, 1977.

%
"Jag vet inte var vi kommer ifrån, Vet inte var vi ska, Och om allt detta skulle ha en anledning, Vi skulle vara den sista att veta. Så låt oss hoppas bara att det är ett förlovat land, Och tills dess, ... Så gott du kan. "
		-- Steppenwolf, "Rock Me Baby"

%
"Hjälp Mr Wizard!"
		-- Tennessee Tuxedo

%
"Den lagstiftare, av alla varelser, beror de flesta lagen trohet. Han av alla män bör bete sig som om lagen tvingade honom. Men det är den universella svaghet för mänskligheten att vad vi är ges att administrera vi nu föreställer vi äger. "
		-- H. G. Wells

%
"Till skillnad från de flesta net.puritans dock känner jag att vad andra samtyckande datorer göra i avskildhet i sina egna telefonförbindelser är deras egen verksamhet. "
		-- John Woods, jfw@eddie.mit.edu

%
"Prata inte med mig om friskrivning! Jag uppfann friskrivning!"
		-- The Censored Hacker

%
"På denna punkt vi vill vara helt klar: socialism har ingenting att göramed utjämning. Socialismen kan inte garantera livsvillkor ochlivsmedel i enlighet med principen "Från var och en efter hansförmåga, åt var och en efter hans behov. "Detta kommer att vara under kommunismen.Socialismen har ett annat kriterium för att fördela sociala förmåner:"Från var och en efter förmåga, åt var och en efter hans arbete." "
		-- Mikhail Gorbachev, _Perestroika_

%
"Cable är inte en lyx, eftersom många områden har dålig TV-mottagning."- Borgmästaren i Tucson, Arizona, 1989[Tydligen är bra TV-mottagning en nödvändighet - åtminstone i Tucson -kl]
		-- Mikhail Gorbachev, _Perestroika_

%
"Alla systemets vägar måste topologiskt och cirkulärt sammankopplade för konceptuellt definitiv lokalt transform, polyhedronal förståelse för uppnås i vår spontana - ergo, mest ekonomiska - geodesiccally strukturerade tankar. "
		-- R. Buckminster Fuller [...and a total nonsequitur as far as I can tell.  -kl]

%
"En sak som de inte berätta om att göra experimentell fysik är att Ibland måste du arbeta under svåra förhållanden ... som ett tillstånd av ren skräck."
		-- W. K. Hartmann

%
"Det är när de säger 2 + 2 = 5 som jag börjar argumentera."
		-- Eric Pepke

%
Jämföra information och kunskap är som att be om fetma av engris är mer eller mindre grön än utsedd slagman regeln. "
		-- David Guaspari

%
"Ingen av våra män är" experter. "Vi har mest tyvärr funnit det nödvändigtatt bli av med en man så snart som han tror sig en expert - eftersom ingennågonsin anser sig expert om han verkligen vet sitt jobb. En man som vetjobb ser så mycket mer att göra än vad han har gjort, att han alltid pressarframåt och aldrig ger upp ett ögonblick av tanke till hur bra och hur effektivthan är. Tänker alltid framåt, tänker alltid att försöka göra mer, ger ensinnestillstånd där ingenting är omöjligt. I det ögonblick man får in i"Expert" state of mind ett stort antal saker blir omöjligt. "
		-- From Henry Ford Sr., "My Life and Work," p. 86 (1922):

%
"NY Times läses av människor som driver landet. The Washington Postläses av människor som tror att de kör landet. National Enquirerläses av människor som tror att Elvis lever och styra landet ... "
		-- Robert J Woodhead (trebor@biar.UUCP)

%
        "..." Eld "spelar ingen roll," jord "och" luft "och" vatten "intemateria. "Jag spelar ingen roll. Inga ord betyder. Men man glömmer verklighetenoch minns ord. Ju fler ord han minns, det smartare att göra sittassistenter uppskattar honom. Han ser på de stora omvandlingen avvärld, men han inte ser dem som de sågs när man såg påverklighet för första gången. Deras namn kommer till sina läppar och han lersom han smakar dem och tänkte att han känner dem i namngivningen. "
		-- Siddartha, _Lord_of_Light_ by Roger Zelazny

%
"Bevattning av landet med havsvatten avsaltas genom fusionskraft är gammal.Det kallas "regn". "
		-- Michael McClary, in alt.fusion

%
"Den dåliga rykte UNIX har fått är helt oförtjänt, som på av människor som inte förstår, som inte har kommit in där och försökte något. "
		-- Jim Joyce, former computer science lecturer at the University of California

%
"Vi forskare, vars tragiska öde har varit att göra de metoder förförintelse alltmer ohyggliga och mer effektiv måste överväga det vår högtidligoch transcendent plikt att göra allt i vår makt för att förhindra dessa vapen frånanvänds för brutal ändamål för vilka de uppfanns. "
		-- Albert Einstein, Bulletin of Atomic Scientists, September 1948

%
"Du kan ha min Unix-system när du bänder det ur mina kalla, döda fingrar."
		-- Cal Keegan

%
Vi kommer mer än gärna göra det en gång Jim visar minsta teckenintresse för fastställande av hans förslag för att ta itu med de tekniskaargument som har * redan * gjorts. De flesta ingenjörer harlärt det finns lite att vinna i finjustera ventiltiderpå en bensindriven förbränningsmotor när kolvarnaoch vevaxel saknas ...
		-- Valdis.Kletnieks@vt.edu on NANOG

%
Det är alltid tråkigt när lopporna lämnar, eftersom det innebär att din hund är död.
		-- Wesley T. Williams

%
