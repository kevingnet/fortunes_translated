BOFH vändning # 1:klockfrekvens

%
BOFH ursäkt # 2:solstormar

%
BOFH ursäkt # 3:elektromagnetisk strålning från satelliten skräp

%
BOFH vändning # 4:statisk från nylon underkläder

%
BOFH ursäkt # 5:statisk från plast räknestickor

%
BOFH vändning # 6:Global uppvärmning

%
BOFH vändning # 7:dålig effektkonditione

%
BOFH vändning # 8:statisk elektricitet

%
BOFH vändning # 9:dopplereffekt

%
BOFH ursäkt # 10:hårdvara stressfrakturer

%
BOFH ursäkt # 11:magnetiska störningar från pengarna / kreditkort

%
BOFH vändning # 12:torra fogar på kabelkontakt

%
BOFH ursäkt # 13:vi väntar på [telefonbolaget] för att åtgärda den linjen

%
BOFH vändning # 14:låter som en Windows-problem, prova att ringa Microsofts support

%
BOFH ursäkt # 15:tillfällig dirigerings anomali

%
BOFH ursäkt # 16:någon var beräkna pi på servern

%
BOFH ursäkt # 17:fett elektroner i ledningarna

%
BOFH ursäkt # 18:överskott överspänningsskydd

%
BOFH ursäkt # 19:flyttalsprocessor spill

%
BOFH ursäkt # 20:dela-med-noll fel

%
BOFH ursäkt # 21:POSIX efterlevnad problem

%
BOFH ursäkt # 22:bildskärmsupplösning för hög

%
BOFH ursäkt # 23:felaktigt orienterad tangentbord

%
BOFH ursäkt # 24:nätverkspaket som reser uppför (använd en bärare duva)

%
BOFH ursäkt # 25:Minskande elektronflöde

%
BOFH ursäkt # 26:första lördagen efter första fullmånen i vinter

%
BOFH ursäkt # 27:radiositet utarmning

%
BOFH ursäkt # 28:CPU radiator bruten

%
BOFH ursäkt # 29:Det fungerar som Wang gjorde, vad är problemet

%
BOFH ursäkt # 30:positron router felfunktion

%
BOFH ursäkt # 31:cellulär telefon interferens

%
BOFH ursäkt # 32:techtonic påkänning

%
BOFH ursäkt # 33:piezoelektrisk störningar

%
BOFH ursäkt # 34:(L) användarfel

%
BOFH ursäkt # 35:fungerar som utformats

%
BOFH ursäkt # 36:dynamisk programvara länkningstabellen skadad

%
BOFH ursäkt # 37:tung allvar fluktuationer, flytta datorn till golvet snabbt

%
BOFH ursäkt # 38:sekreterare inkopplad hårtork till UPS

%
BOFH ursäkt # 39:terroristverksamhet

%
BOFH ursäkt # 40:inte tillräckligt med minne, gå och hämta systemuppgradering

%
BOFH ursäkt # 41:avbrotts konfigurationsfel

%
BOFH ursäkt # 42:spagetti kabel orsakar paket misslyckande

%
BOFH ursäkt # 43:boss glömt systemlösenord

%
BOFH ursäkt # 44:helgdag - systemet rörelsekrediter inte laddas

%
BOFH ursäkt # 45:virus attack, loser ansvarig

%
BOFH ursäkt # 46:avloppsvatten tank spill på dator

%
BOFH ursäkt # 47:Komplett Transient Lockout

%
BOFH ursäkt # 48:dålig eter i kablarna

%
BOFH ursäkt # 49:bogon utsläpp

%
BOFH ursäkt # 50:Förändring i jordens rotationshastighet

%
BOFH ursäkt # 51:Kosmisk strålning partiklar kraschade igenom hårddisken tallrik

%
BOFH ursäkt # 52:Lukt från ohygieniska vaktmästeri personal havererade bandhuvudena

%
BOFH ursäkt # 53:Lilla hamstern i löphjul hade krans; väntar på byte som skall Fedexed från Wyoming

%
BOFH ursäkt # 54:Onda hundar hypnotiserade nattskift

%
BOFH ursäkt # 55:Plumber misstog routing panel för dekorativa väggfäste

%
BOFH ursäkt # 56:Elektriker gjorde popcorn i strömförsörjningen

%
BOFH ursäkt # 57:Vårdare stal root-lösenordet

%
BOFH ursäkt # 58:systemfel högtrycks

%
BOFH ursäkt # 59:misslyckade försök, systembehov omgjorda

%
BOFH ursäkt # 60:Systemet har återkallats

%
BOFH ursäkt # 61:inte godkänts av FCC

%
BOFH ursäkt # 62:behöver svepa systemet i aluminiumfolie för att åtgärda problemet

%
BOFH ursäkt # 63:inte ordentligt jordad, vänligen begrava dator

%
BOFH ursäkt # 64:CPU behöver kalibreras

%
BOFH ursäkt # 65:systemet behöver startas om

%
BOFH ursäkt # 66:bitbucket overflow

%
BOFH ursäkt # 67:avkoda kod behövs från mjukvaruföretag

%
BOFH ursäkt # 68:endast tillgänglig på ett behov av att veta grunden

%
BOFH ursäkt # 69:knut i kablar orsakade dataströmmen att bli vridna och snodd

%
BOFH ursäkt # 70:häckande kackerlackor sluten ut eter kabel

%
BOFH ursäkt # 71:Filsystemet är fullt av det

%
BOFH ursäkt # 72:Satan gjorde det

%
BOFH ursäkt # 73:Demoner gjorde det

%
BOFH ursäkt # 74:Du är slut på minne

%
BOFH ursäkt # 75:Det finns inte några problem

%
BOFH ursäkt # 76:Unoptimized hårddisk

%
BOFH ursäkt # 77:Stavfel i koden

%
BOFH ursäkt # 78:Ja, ja, det som kallas ett designbegränsning

%
BOFH ursäkt # 79:Titta, kompis: Windows 3.1 är en allmän skyddsfel.

%
BOFH ursäkt # 80:Det är en stor dator du har där; har du funderat på hur det skulle fungera som en BSD maskin?

%
BOFH ursäkt # 81:Ursäkta mig, jag har till kretsen en växelströmsledning genom mitt huvud att få denna databas arbets.

%
BOFH ursäkt # 82:Ja, yo mama klänningar du roliga och du behöver en mus för att radera filer.

%
BOFH ursäkt # 83:Stödpersonal bakfull, skicka aspirin och komma tillbaka senare.

%
BOFH ursäkt # 84:Någon står på Ethernet-kabel, vilket orsakar en knut i kabeln

%
BOFH ursäkt # 85:Windows 95 papperslösa "funktion"

%
BOFH ursäkt # 86:Runt paket

%
BOFH ursäkt # 87:Lösenordet är för komplex för att dekryptera

%
BOFH ursäkt # 88:Boss 'unge fucked up maskinen

%
BOFH ursäkt # 89:Elektromagnetisk energiförlust

%
BOFH ursäkt # 90:Budgetnedskärningar

%
BOFH ursäkt # 91:Mus tuggas genom strömkabel

%
BOFH ursäkt # 92:Unken fil handtag (nästa gång använda Tupperware (tm)!)

%
BOFH ursäkt # 93:Har ännu inte genomförts

%
BOFH ursäkt # 94:internet strömavbrott

%
BOFH ursäkt # 95:Pentium Fdiv Bugg

%
BOFH ursäkt # 96:Leverantör inte längre stöder produkten

%
BOFH ursäkt # 97:Små djur kamikaze attack på nätaggregat

%
BOFH ursäkt # 98:Säljaren sätta bugg där.

%
BOFH ursäkt # 99:SIMM överhörning.

%
BOFH ursäkt # 100:IRQ dropout

%
BOFH ursäkt # 101:hopfällda Backbone

%
BOFH ursäkt # 102:Power Company testa nya spänningsspiken (skapande) utrustning

%
BOFH ursäkt # 103:operatörer i strejk på grund av brutna kaffebryggare

%
BOFH ursäkt # 104:backup band över med kopia av System Manager favorit CD

%
BOFH ursäkt # 105:UPS avbröt serverns makt

%
BOFH ursäkt # 106:Elektrikern visste inte vad den gula kabeln var så han ryckte ethernet ut.

%
BOFH ursäkt # 107:Tangentbordet är inte ansluten

%
BOFH ursäkt # 108:Luftkonditioneringen vattenledningen spruckit över maskinrummet

%
BOFH ursäkt # 109:Den el transformatorstation på parkeringen sprängdes.

%
BOFH ursäkt # 110:Rolling Stones konsert på vägen orsakade en brun ut

%
BOFH ursäkt # 111:Försäljaren körde över CPU-kortet.

%
BOFH ursäkt # 112:Bildskärmen är ansluten till den seriella porten

%
BOFH ursäkt # 113:Root namnservrar är ur synk

%
BOFH ursäkt # 114:elektromagnetiska pulser från Franska ovan jord nuke testning.

%
BOFH ursäkt # 115:tangentbordets mellanslagstangenten genererar falska tangentkoder.

%
BOFH ursäkt # 116:de verkliga ttys blev pseudo ttys och vice versa.

%
BOFH ursäkt # 117:skrivaren tänker dess en router.

%
BOFH ursäkt # 118:routern tänker dess en skrivare.

%
BOFH ursäkt # 119:onda hackare från Serbien.

%
BOFH ursäkt # 120:vi bara bytt till FDDI.

%
BOFH ursäkt # 121:halon systemet gick och dödade operatörerna.

%
BOFH ursäkt # 122:eftersom Bill Gates är ett Jehovas vittne och så ingenting kan arbeta på St Swithin dag.

%
BOFH ursäkt # 123:användaren att datorförhållande för hög.

%
BOFH ursäkt # 124:användaren att datorn ranson för låg.

%
BOFH ursäkt # 125:vi bara bytt till Sprint.

%
BOFH ursäkt # 126:Det har Intel Inside

%
BOFH ursäkt # 127:Klibbiga bitar på disk.

%
BOFH ursäkt # 128:Power Company har EMP problem med sin reaktor

%
BOFH ursäkt # 129:Ringen behöver en annan token

%
BOFH ursäkt # 130:ny ledning

%
BOFH ursäkt # 131:telnet: Kan inte ansluta till fjärrvärden: Connection refused

%
BOFH ursäkt # 132:SCSI Chain overterminated

%
BOFH ursäkt # 133:Det är inte inkopplad.

%
BOFH ursäkt # 134:på grund av nätverks eftersläpning på grund av för många personer som spelar deathmatch

%
BOFH ursäkt # 135:Du sätter skivan i upp och ned.

%
BOFH ursäkt # 136:Demoner löst i systemet.

%
BOFH ursäkt # 137:Användar delade ut pornografi på servern; Systemet beslagtagits av FBI.

%
BOFH ursäkt # 138:BNC (hjärna inte ansluten)

%
BOFH ursäkt # 139:UBNC (användar hjärnan inte ansluten)

%
BOFH ursäkt # 140:LBNC (loser hjärnan inte ansluten)

%
BOFH ursäkt # 141:diskar snurrar bakåt - växla halvklotet bygeln.

%
BOFH ursäkt # 142:nya killen korskopplade telefonlinjer med växelströmsbussen.

%
BOFH ursäkt # 143:var tvungen att använda hammare för att frigöra fastnat hårddisk huvuden.

%
BOFH ursäkt # 144:Alltför få computrons tillgängliga.

%
BOFH ursäkt # 145:Punktering på herrgårdsvagn med band. ( "Underskatta aldrig bandbredden för en stationsvagn full av band slunga på motorvägen" Andrew S. Tannenbaum)

%
BOFH ursäkt # 146:Kommunikationssatellit som används av militären för star wars.

%
BOFH ursäkt # 147:Party-bugg i Aloha-protokollet.

%
BOFH ursäkt # 148:Sätt mynt för nytt spel

%
BOFH ursäkt # 149:Dagg på telefonlinjer.

%
BOFH vändning # 150:ARCserve kraschade servern igen.

%
BOFH ursäkt # 151:Någon behövde powerstrip, så de drog växeln kontakten.

%
BOFH ursäkt # 152:Min hästsvans träffade på / av-knapp på grenuttag.

%
BOFH ursäkt # 153:Stort att little endian konvertering fel

%
BOFH ursäkt # 154:Du kan ställa ett filsystem, men du kan inte ställa in en fisk (från de flesta tunefs manualsidor)

%
BOFH ursäkt # 155:dum terminal

%
BOFH ursäkt # 156:Zombie processer spöka datorn

%
BOFH ursäkt # 157:Felaktig tidssynkronisering

%
BOFH ursäkt # 158:nedlagda processer

%
BOFH ursäkt # 159:envisa processer

%
BOFH ursäkt # 160:icke-redundant fläktfel

%
BOFH ursäkt # 161:övervaka VLF läckage

%
BOFH ursäkt # 162:buggar i RAID

%
BOFH ursäkt # 163:nej "någon" tangent på tangentbordet

%
BOFH ursäkt # 164:rotröta

%
BOFH ursäkt # 165:backbone skolios

%
BOFH ursäkt # 166:/ Pub / lunch

%
BOFH ursäkt # 167:drivna kollisioner och inte tillräckligt paket ambulanser

%
BOFH ursäkt # 168:le0: ingen bärvåg: transceiver kabel problem?

%
BOFH ursäkt # 169:sända paket på fel frekvens

%
BOFH ursäkt # 170:popper inte behandla jumbo kärna

%
BOFH ursäkt # 171:OBSERVERA: Alloc: / dev / null: filsystem fullt

%
BOFH ursäkt # 172:pseudo-användare på en pseudo-terminal

%
BOFH ursäkt # 173:Rekursiv genomgång av loopback monteringspunkter

%
BOFH ursäkt # 174:backbone justering

%
BOFH ursäkt # 175:OS bytte till disk

%
BOFH ursäkt # 176:ångor från avdunstande klibbig-notera lim

%
BOFH ursäkt # 177:sticktion

%
BOFH ursäkt # 178:korta benet på processbord

%
BOFH ursäkt # 179:multicast på trasiga paketen

%
BOFH ursäkt # 180:eter läcka

%
BOFH ursäkt # 181:Atilla hubben

%
BOFH ursäkt # 182:endotermisk omkalibrering

%
BOFH ursäkt # 183:filsystem inte tillräckligt stor för Jumbo Kernel Patch

%
BOFH ursäkt # 184:slinga finns i en slinga i redundant loopback

%
BOFH ursäkt # 185:Systemet konsumerade alla papper för personsökning

%
BOFH ursäkt # 186:åtkomst nekad

%
BOFH ursäkt # 187:Omformatering Page. Vänta...

%
BOFH ursäkt # 188:..disk eller processorn är i brand.

%
BOFH ursäkt # 189:SCSI är för bred.

%
BOFH ursäkt # 190:Proprietary Information.

%
BOFH ursäkt # 191:Skriv bara "mv * / dev / null".

%
BOFH ursäkt # 192:skenande katt på systemet.

%
BOFH ursäkt # 193:Har du betala nya Support Fee?

%
BOFH ursäkt # 194:Vi stöder bara en 1200 bps-anslutning.

%
BOFH ursäkt # 195:Vi stöder bara en 28000 bps anslutning.

%
BOFH ursäkt # 196:Mig inga internet, bara vaktmästare, jag bara vax golv.

%
BOFH ursäkt # 197:Jag är ledsen en Pentium kommer inte att göra, behöver du en SGI att ansluta med oss.

%
BOFH ursäkt # 198:Post-it-lapp Slam läckt in i monitorn.

%
BOFH ursäkt # 199:lockarna i tangentbordet sladd förlorar el.

%
BOFH ursäkt # 200:Monitorn behöver en annan låda av pixlar.

%
BOFH ursäkt # 201:RPC_PMAP_FAILURE

%
BOFH ursäkt # 202:kernel panic: skriva-only-minne (/ dev / wom0) kapacitet överskrids.

%
BOFH ursäkt # 203:Skriv-only-minne delsystem för långsam för denna maskin. Kontakta din lokala återförsäljare.

%
BOFH ursäkt # 204:Bara plocka upp telefonen och ge modem ansluta ljud. "Ja du sa att vi skulle få fler linjer så att vi inte har linjer."

%
BOFH ursäkt # 205:Kvantdynamik påverkar transistorerna

%
BOFH ursäkt # 206:Polisen undersöker alla internetpaket i sökandet efter en knarknettohandlare

%
BOFH ursäkt # 207:Vi är för närvarande försöker ett nytt koncept för att använda en levande mus. Tyvärr har en ännu överleva som ansluten till datorn ..... tänk med oss.

%
BOFH ursäkt # 208:Din e-post dirigeras genom Tyskland ... och de är censurera oss.

%
BOFH ursäkt # 209:Endast personer med namn som börjar med "A" får post denna vecka (a la Microsoft)

%
BOFH ursäkt # 210:Vi betalade inte Internet räkningen och det har varit avskuren.

%
BOFH ursäkt # 211:Blixtnedslag.

%
BOFH ursäkt # 212:Naturligtvis är det inte fungerar. Vi har utfört en mjukvaruuppgradering.

%
BOFH ursäkt # 213:Ändra språk till finska.

%
BOFH ursäkt # 214:Lysrör genererar negativa joner. Om stänga av dem inte fungerar, ta ut dem och sätta aluminiumfolie på ändarna.

%
BOFH ursäkt # 215:Hög kärnteknisk verksamhet i ditt område.

%
BOFH ursäkt # 216:Vad kontor är du i? Åh, att en. Visste du att byggnaden byggdes över universitet första kärnforskningsanläggning? Och wow, är inte du den lycklige, kontoret är rätt över där kärnan är begravd!

%
BOFH ursäkt # 217:MGS slut på gas.

%
BOFH ursäkt # 218:UPS har inte en batteribackup.

%
BOFH ursäkt # 219:Recursivity. Ring tillbaka om det händer igen.

%
BOFH ursäkt # 220:Någon trodde den stora röda knappen var en strömbrytare.

%
BOFH ursäkt # 221:Stordatorn behöver vila. Det börjar bli gammal, du vet.

%
BOFH ursäkt # 222:Jag är inte säker. Försök att ringa Internet huvudkontor - det är i boken.

%
BOFH ursäkt # 223:Linjerna är alla upptagna (busied ut, det vill säga - varför låt dem till att börja med).

%
BOFH ursäkt # 224:9 januari 16:41:27 Huber SU: "su root" lyckats för .... på / dev / pts / 1

%
BOFH ursäkt # 225:Det är de dator människor i X {staden av världs}. De håller upp fyllning saker.

%
BOFH ursäkt # 226:En star wars satellit misstag sprängde WAN.

%
BOFH vändning # 227:Allvarligt fel rakt framför skärmen

%
BOFH ursäkt # 228:Denna funktion är för närvarande inte stöds, men Bill Gates försäkrar oss att det kommer att finnas med i nästa uppgradering.

%
BOFH ursäkt # 229:fel polaritet neutron flöde

%
BOFH ursäkt # 230:Lusers inlärningskurva verkar vara fraktal

%
BOFH ursäkt # 231:Vi var tvungna att stänga av tjänsten att följa CDA Bill.

%
BOFH ursäkt # 232:Jonisering från luftkonditionerings

%
BOFH ursäkt # 233:TCP / IP UDP larmgränsen är satt för lågt.

%
BOFH ursäkt # 234:Någon sänder pygmé paket och routern inte vet hur man handskas med dem.

%
BOFH ursäkt # 235:Den nya frame relay nätverk har inte bäddas ner programvaran slingan sändaren ännu.

%
BOFH ursäkt # 236:Fanout släppa spänningen för mycket, försök skära några av dessa små spår

%
BOFH ursäkt # 237:Platta spänning för lågt på demodulator rör

%
BOFH ursäkt # 238:Du gjorde wha ... oh _dear _....

%
BOFH ursäkt # 239:Centralprocessorer kullager omförpackade

%
BOFH ursäkt # 240:Alltför många små stift på CPU förvirrande det, böja fram och tillbaka tills 10-20% är snyggt bort. Gör _inte_ lämna metallbitar synlig!

%
BOFH ursäkt # 241:_Rosin_ Kärna löda? Men...

%
BOFH ursäkt # 242:Software använder amerikanska mått, men OS är i metriska ...

%
BOFH ursäkt # 243:Datorn fleetly, mus och alla.

%
BOFH ursäkt # 244:Din katt försökte äta musen.

%
BOFH ursäkt # 245:Borg försökte assimilera datorn. Motstånd är meningslöst.

%
BOFH ursäkt # 246:Det måste ha varit åskväder hade vi (igår) (förra veckan) (förra månaden)

%
BOFH ursäkt # 247:På grund av federala problem budget vi har varit tvungna att skära ner på antalet användare som kan få tillgång till systemet på en gång. (Det vill säga ingen tillåten ....)

%
BOFH ursäkt # 248:För mycket strålning som kommer från marken.

%
BOFH ursäkt # 249:Tyvärr har vi slut på bitar / bytes / vad som helst. Oroa dig inte, kommer nästa leverans komma nästa vecka.

%
BOFH ursäkt # 250:Program belastning för tung för processorn att lyfta.

%
BOFH ursäkt # 251:Processer som körs långsamt på grund av svag strömförsörjning

%
BOFH ursäkt # 252:Vår ISP har {omkopplings, routing, SMD, frame relay} problem

%
BOFH ursäkt # 253:Vi har slut på licenser

%
BOFH ursäkt # 254:Störningar från månens strålning

%
BOFH ursäkt # 255:Stående rum bara på bussen.

%
BOFH ursäkt # 256:Du måste installera ett RTFM gränssnitt.

%
BOFH ursäkt # 257:Det skulle bero på att programmet inte fungerar.

%
BOFH ursäkt # 258:Det är lätt att fixa, men jag kan inte bli störd.

%
BOFH ursäkt # 259:Någon tie fångas i skrivaren, och om något annat blir tryckt, kommer han att vara i det också.

%
BOFH ursäkt # 260:Vi uppgraderar / dev / null

%
BOFH ursäkt # 261:Usenet nyheten är inaktuell

%
BOFH ursäkt # 262:Vår POP server kidnappades av en vessla.

%
BOFH ursäkt # 263:Det har fastnat på webben.

%
BOFH ursäkt # 264:Modemet inte talar engelska.

%
BOFH ursäkt # 265:Musen rymt.

%
BOFH ursäkt # 266:Alla paketen är tomma.

%
BOFH ursäkt # 267:UPS-enheten är i strejk.

%
BOFH ursäkt # 268:Neutrino överbelastning på namnservern

%
BOFH ursäkt # 269:Smältande hårddiskar

%
BOFH ursäkt # 270:Någon har trasslat till kärnan pekare

%
BOFH ursäkt # 271:Kärnan licens har gått ut

%
BOFH ursäkt # 272:Netscape har kraschat

%
BOFH ursäkt # 273:Sladden hoppade över och slå på strömbrytaren.

%
BOFH ursäkt # 274:Det var OK innan du rörde vid den.

%
BOFH ursäkt # 275:bitars röta

%
BOFH ursäkt # 276:US Postal Service

%
BOFH ursäkt # 277:Din Flux Kondensator har gått dåligt.

%
BOFH ursäkt # 278:De Dilithium Kristaller måste roteras.

%
BOFH ursäkt # 279:Den statiska elektricitet routing handlar upp ...

%
BOFH ursäkt # 280:Traceroute säger att det finns en dirigeringsproblem i huvudkedjan. Det är inte vårt problem.

%
BOFH ursäkt # 281:Co-locator kan inte verifiera frame-relay inkörsport till ISDN-servern.

%
BOFH ursäkt # 282:Hög höjd kondens från U.S.A.F prototyp flygplan har förorenat den primära nätmask. Stäng av datorn för 9 dagar för att undvika att skada den.

%
BOFH ursäkt # 283:Gräsklippare blad i din fan behöver vässa

%
BOFH ursäkt # 284:Elektroner på en bender

%
BOFH ursäkt # 285:Telekommunikation uppgraderar.

%
BOFH ursäkt # 286:Telekommunikation är nedgradering.

%
BOFH ursäkt # 287:Telekommunikation nedväxling.

%
BOFH ursäkt # 288:Hårddisk sova. Låt den vakna upp på egen hand ...

%
BOFH ursäkt # 289:Interferens mellan tangentbordet och stolen.

%
BOFH ursäkt # 290:Processorn har skiftat, och blir decentraliserat.

%
BOFH ursäkt # 291:På grund av CDA, vi inte längre har en root-kontot.

%
BOFH ursäkt # 292:Vi har slut på kopplingston och vi och väntar på telefonbolaget för att leverera en annan flaska.

%
BOFH ursäkt # 293:Du måste ha slå fel på valfri tangent.

%
BOFH ursäkt # 294:PCMCIA slavdrivare

%
BOFH ursäkt # 295:Token föll ut ur ringen. Ring oss när du hittar den.

%
BOFH ursäkt # 296:Hårdvaran buss behöver en ny token.

%
BOFH ursäkt # 297:Alltför många avbrott

%
BOFH ursäkt # 298:Inte tillräckligt avbrott

%
BOFH ursäkt # 299:Data på hårddisken är ur balans.

%
BOFH ursäkt # 300:Digital Manipulator överskrider hastighetsparametrar

%
BOFH ursäkt # 301:verkar vara en långsam / Narrow SCSI-0-gränssnitt problem

%
BOFH ursäkt # 302:mikro Riemannsk krökta rymd fel i skrivskyddat filsystem

%
BOFH ursäkt # 303:fraktal strålning fastnar ryggraden

%
BOFH ursäkt # 304:routing problem på neuronnätet

%
BOFH ursäkt # 305:IRQ-problem med Un avbrotts-Power-Supply

%
BOFH ursäkt # 306:CPU-vinkel har justeras på grund av vibrationer som kommer från närliggande väg

%
BOFH ursäkt # 307:utsläpp från GSM-telefoner

%
BOFH ursäkt # 308:CD-ROM-server behöver kalibreras

%
BOFH ursäkt # 309:Brandväggen behöver kylning

%
BOFH ursäkt # 310:asynkron inod misslyckande

%
BOFH ursäkt # 311:gående bussprotokoll kränkning

%
BOFH ursäkt # 312:inkompatibla bit registrerings operatörer

%
BOFH ursäkt # 313:din process är inte ISO 9000-kompatibel

%
BOFH ursäkt # 314:Du måste uppgradera din VESA lokalbuss till en Masterlokalbuss.

%
BOFH ursäkt # 315:Den senaste tidens spridning av kärnvapenprov

%
BOFH ursäkt # 316:Älvor i strejk. (Varför de kallar EMAG Elf Magi)

%
BOFH ursäkt # 317:Internet översteg Luser nivå, vänta tills en loser loggar ut innan du försöker logga in igen.

%
BOFH ursäkt # 318:Din e-postadress är nu levereras av USPS.

%
BOFH ursäkt # 319:Datorn har inte återvänder alla bitar det blir från Internet.

%
BOFH ursäkt # 320:Du har blivit smittad av teleskop Hubble-viruset.

%
BOFH ursäkt # 321:Planerad global CPU strömavbrott

%
BOFH ursäkt # 322:Din Pentium har en värmeproblem - prova kylning med iskallt vatten (Stäng inte av datorn, vill du inte att kyla ner Pentium Chip när han inte fungerar, eller hur?).

%
BOFH ursäkt # 323:Din processor har bearbetat för många instruktioner. Stäng av den omedelbart, inte skriva några kommandon !!

%
BOFH ursäkt # 324:Dina paket var uppätna av terminatorn

%
BOFH ursäkt # 325:Din processor utvecklar inte tillräckligt med värme.

%
BOFH ursäkt # 326:Vi behöver en behörig elektriker för att ersätta glödlampor i datasalen.

%
BOFH ursäkt # 327:POP-servern är ur koks

%
BOFH ursäkt # 328:Fiberoptik orsakade gas huvud läcka

%
BOFH ursäkt # 329:Server deprimerad, behöver Prozac

%
BOFH ursäkt # 330:quantum decoherence

%
BOFH ursäkt # 331:dessa jävla fladdermöss!

%
BOFH ursäkt # 332:suboptimal dirigering erfarenhet

%
BOFH ursäkt # 333:En rörmokare behövs är nätverks avloppet tilltäppta

%
BOFH ursäkt # 334:50% av handboken är i pdf Readme-filen

%
BOFH ursäkt # 335:AA batterier i Väggklocka sänder magnetisk störning

%
BOFH ursäkt # 336:xy axel i styrkulan samordnas med sommarsolståndet

%
BOFH ursäkt # 337:butan tändaren bringar pincushioning

%
BOFH ursäkt # 338:gamla bläckpatroner härrör barium baserade rök

%
BOFH ursäkt # 339:chef i ledningskanalen

%
BOFH ursäkt # 340:Väl fixa det i nästa (uppgradering, uppdatera patch release, service pack).

%
BOFH ursäkt # 341:HTTPD Fel 666: BOFH var här

%
BOFH ursäkt # 342:HTTPD Fel 4004: mycket gamla Intel CPU - otillräcklig processorkraft

%
BOFH ursäkt # 343:ATM styrelse har slut på 10 pundsedlar. Vi har en piska runt för att fylla på den, till vård bidra?

%
BOFH ursäkt # 344:Nätverksfel - ring NBC

%
BOFH ursäkt # 345:Att manuellt spåra satelliten.

%
BOFH ursäkt # 346:Din / vår dator (s) hade drabbats av en minnesläcka, och vi väntar på att de ska fyllas på.

%
BOFH ursäkt # 347:Gummibandet bröt

%
BOFH ursäkt # 348:Vi är på Token Ring, och det ser ut som token fick loss.

%
BOFH ursäkt # 349:Stray alfapartiklar från minnet förpackning orsakade Hard minnesfel på servern.

%
BOFH ursäkt # 350:paradigmskifte ... utan en koppling

%
BOFH ursäkt # 351:PEBKAC (Problem finns mellan tangentbord och ordförande)

%
BOFH ursäkt # 352:Kablarna är inte samma längd.

%
BOFH ursäkt # 353:Second-systemet effekt.

%
BOFH ursäkt # 354:Tuggummi på / dev / sd3c

%
BOFH ursäkt # 355:Tristess i kärnan.

%
BOFH ursäkt # 356:de demoner! de demoner! de fruktansvärda demoner!

%
BOFH ursäkt # 357:Jag vill gärna hjälpa dig - det är bara att chefen inte kommer att låta mig i närheten av datorn.

%
BOFH ursäkt # 358:slås av Good Times-virus

%
BOFH ursäkt # 359:DU ETT I / O-FEL -> inkompetent operatörsfel

%
BOFH ursäkt # 360:Din paritetskontroll är övertrasserat och du är ute cache.

%
BOFH ursäkt # 361:Kommunistiska revolutionärer tar över serverrummet och krävande alla datorer i huset eller de skjuter sysadmin. Dåliga vilseledda dårar.

%
BOFH ursäkt # 362:Plasmaledningsbrott

%
BOFH ursäkt # 363:Av korten på enhet D:

%
BOFH ursäkt # 364:Sand loppor äter Internet kablar

%
BOFH ursäkt # 365:parallella processorer löper vinkelrätt idag

%
BOFH ursäkt # 366:ATM-cell har ingen roaming-funktionen aktiverad, kan bärbara datorer inte ansluta

%
BOFH ursäkt # 367:Webmasters kidnappad av onda kult.

%
BOFH ursäkt # 368:Underlåtenhet att justera för sommartid.

%
BOFH ursäkt # 369:Virus som överförs från datorn till systemadministratörer.

%
BOFH ursäkt # 370:Virus på grund av datorer som har det osäkra könet.

%
BOFH ursäkt # 371:Felaktigt konfigurerade statiska vägar på corerouters.

%
BOFH ursäkt # 372:Tvingad att stödja NT-servrar; sysadmins sluta.

%
BOFH ursäkt # 373:Misstänkta pekare skadad virtuell maskin

%
BOFH ursäkt # 374:Det är InterNIC fel.

%
BOFH ursäkt # 375:Rotnamnsservrar skadad.

%
BOFH ursäkt # 376:budgetnedskärningar tvingade oss att sälja alla strömkablar för servrarna.

%
BOFH ursäkt # 377:Någon fast de partvinnade ledningarna till telefonsvararen.

%
BOFH ursäkt # 378:Operatörer som dödats av år 2000 bugg bita.

%
BOFH ursäkt # 379:Vi har plockat COBOL som språkvalet.

%
BOFH ursäkt # 380:Operatörer dödades när jättehög med backup band föll.

%
BOFH ursäkt # 381:Robotic band växlare misstog operatörens oavgjort för en backup band.

%
BOFH ursäkt # 382:Någon rökning i datasalen och kvitta halonsystemen.

%
BOFH ursäkt # 383:Din processor har tagit en tur till Heaven Gate på UFO bakom Hale-Bopp komet.

%
BOFH ursäkt # 384:Det är ett ID-10-T-fel

%
BOFH ursäkt # 385:Dyslektiker skriva om hosts på servrar

%
BOFH ursäkt # 386:Internet genomsöks efter virus.

%
BOFH ursäkt # 387:Datorns fackliga avtal är inställd på att löpa ut vid midnatt.

%
BOFH ursäkt # 388:Dålig användar karma.

%
BOFH ursäkt # 389:/ Dev / ledtråd var kopplat till / dev / null

%
BOFH ursäkt # 390:Ökad solfläcksaktiviteten.

%
BOFH ursäkt # 391:Vi har redan skickat runt ett meddelande om detta.

%
BOFH ursäkt # 392:Det är unionens regler. Det finns inget vi kan göra åt det. Förlåt.

%
BOFH ursäkt # 393:Störningar från Van Allen Belt.

%
BOFH ursäkt # 394:Jupiter är i linje med Mars.

%
BOFH ursäkt # 395:Redundanta ACL.

%
BOFH ursäkt # 396:E-postserver drabbats av UniSpammer.

%
BOFH ursäkt # 397:T-1: s överbelastade på grund av porr trafik till nyhetsservern.

%
BOFH ursäkt # 398:Data för intranät fick dirigeras genom extranät och landade på internet.

%
BOFH ursäkt # 399:Vi är en 100% Microsoft Shop.

%
BOFH ursäkt # 400:Vi är Microsoft. Vad du upplever är inte ett problem; det är ett papperslösa funktionen.

%
BOFH ursäkt # 401:Säljare sålt en produkt som vi inte erbjuda.

%
BOFH ursäkt # 402:Sekreterare skickade kedjebrev till alla 5000 anställda.

%
BOFH ursäkt # 403:Sysadmin hörde inte sökare gå av på grund av hög musik från bar-rums högtalare.

%
BOFH ursäkt # 404:Sysadmin misstag förstörde personsökare med en stor hammare.

%
BOFH ursäkt # 405:Sysadmins otillgängliga eftersom de är i ett möte att tala om varför de inte är tillgängliga så mycket.

%
BOFH ursäkt # 406:Bad kafeteriamat landade alla systemadministratörer på sjukhuset.

%
BOFH ursäkt # 407:Route fladdrande på NAP.

%
BOFH ursäkt # 408:Datorer under vatten på grund av SYN översvämningar.

%
BOFH ursäkt # 409:Vulcan-död-grepp ping har tillämpats.

%
BOFH ursäkt # 410:Elektriska ledningar i maskinrummet smälter.

%
BOFH ursäkt # 411:Trafikstockning på de elektroniska motorvägarna.

%
BOFH ursäkt # 412:Radiell Telemetry Infiltration

%
BOFH ursäkt # 413:Ko-tipp tippas en ko på servern.

%
BOFH ursäkt # 414:Tachyon utsläpp överbelastning av systemet

%
BOFH ursäkt # 415:Underhållsfönster bruten

%
BOFH ursäkt # 416:Vi är ute spår på servern

%
BOFH ursäkt # 417:Datorrum flyttas. Våra system är nere för helgen.

%
BOFH ursäkt # 418:Sysadmins upptagen slåss SPAM.

%
BOFH ursäkt # 419:Upprepade omstarter av systemet misslyckats med att lösa problemet

%
BOFH ursäkt # 420:Funktionen var inte beta testats

%
BOFH ursäkt # 421:Domänkontrollant svarar inte

%
BOFH ursäkt # 422:Någon annan stal din IP-adress, ringa Internet detektiver!

%
BOFH ursäkt # 423:Det är inte RFC-822-kompatibel.

%
BOFH ursäkt # 424:Åtgärden misslyckades eftersom: det finns inget meddelande för detta fel (# 1014)

%
BOFH ursäkt # 425:stoppbit fått

%
BOFH ursäkt # 426:behövs internet för att fånga etherbunny

%
BOFH ursäkt # 427:nätverk ner, IP-paket som levereras via UPS

%
BOFH ursäkt # 428:Firmware uppdatering i kaffemaskinen

%
BOFH ursäkt # 429:temporal anomali

%
BOFH ursäkt # 430:Musen har out-of-ost-error

%
BOFH ursäkt # 431:Borg implantat misslyckas

%
BOFH ursäkt # 432:Borg naniter har angripna servern

%
BOFH ursäkt # 433:error: en dålig användar finns framför skärmen

%
BOFH ursäkt # 434:Vänligen ange vilken typ av teknisk nödsituation

%
BOFH ursäkt # 435:Internet stängdes på grund av underhålls

%
BOFH ursäkt # 436:Daemon rymt från pentagram

%
BOFH ursäkt # 437:cirklarna i majs skal

%
BOFH ursäkt # 438:biten har lossnat

%
BOFH ursäkt # 439:Hot Java har gått kallt

%
BOFH ursäkt # 440:Cache miss - ta bättre sikta nästa gång

%
BOFH ursäkt # 441:Hashtabell har woodworm

%
BOFH ursäkt # 442:Trojansk häst har slut på hö

%
BOFH ursäkt # 443:Zombie processer detekteras, maskin hemsöks.

%
BOFH ursäkt # 444:overflow fel i / dev / null

%
BOFH ursäkt # 445:Webbläsare cookie är skadad - någon har varit knapra på det.

%
BOFH ursäkt # 446:Mailer-daemon är upptagen bränna ditt budskap i helvetet.

%
BOFH ursäkt # 447:Enligt Microsoft är det avsiktligt

%
BOFH ursäkt # 448:vi måste uppgraderas till VII

%
BOFH ursäkt # 449:greenpeace free'd de mallocs

%
BOFH ursäkt # 450:Terrorister kraschade ett flygplan i serverrummet, måste ta bort / bin / laden. (Rm -rf / bin / laden)

%
BOFH ursäkt # 451:astropneumatic oscillationer i vattenkylning

%
BOFH ursäkt # 452:Någon körde operativsystemet genom en stavningskontroll.

%
BOFH ursäkt # 453:Spider angrepp i varma fall delar

%
