En KOD för etiskt beteende för patienter:1. INTE FÖRVÄNTA din läkare för att DELA obehaget.Engagemang med patientens lidande kan få honom att förloravärdefulla vetenskaplig objektivitet.2. sig glada hela tiden.Läkaren leder en upptagen och försöker liv och kräver allamildhet och trygghet han kan få.3. Försök att drabbas av sjukdom som du behandlas.Kom ihåg att din läkare har en professionell rykte att upprätthålla.
		-- Dave Barry, "Stay Fit & Healthy Until You're Dead"

%
En KOD för etiskt beteende för patienter:4. inte klaga om behandlingen underlåter att göra lättnad.Du måste tro att din läkare har uppnått en djup insikt isanna natur din sjukdom, som överskrider alla enbart permanentfunktionshinder du har upplevt.5. frågar aldrig din läkare förklara vad han gör eller varför han gör det.Det är förmätet att tro att sådana djupa frågor kan varaförklaras i termer som du skulle förstå.6. SKICKA nya EXPERIMANTAL BEHANDLING lättare.Även om operationen inte kan gynna dig direkt, den resulterandeuppsats kommer säkert att vara av stort intresse.
		-- Dave Barry, "Stay Fit & Healthy Until You're Dead"

%
En KOD för etiskt beteende för patienter:7. betala din medicinska räkningar snabbt och villigt.Du bör överväga det som ett privilegium att bidra, men blygsamt,till välbefinnande av läkare och andra humanister.8. inte lider av sjukdomar som du inte har råd.Det är ren arrogans att ingå avtal sjukdomar som ligger utanför ditt sätt.9. REVEAL aldrig någon av de brister som uppdagats i KURSEN   AV BEHANDLING av din läkare.Patient och läkare relation är en privilegierad en, och du har enheliga plikt att skydda honom från exponering.10. DIE aldrig under i läkarens NÄRVARO eller under hans direkt vård.Detta kommer bara att orsaka honom onödigt besvär och förlägenhet.
		-- Dave Barry, "Stay Fit & Healthy Until You're Dead"

%
En upprörd patienten ringde henne läkarmottagning. "Var det sant", kvinnanfrågade, "att medicinen läkaren hade ordinerats var för restenav sitt liv? "Hon fick veta att det var. Det fanns bara ett ögonblick av tystnad innankvinnan fortsatte tappert vidare. "Jo, jag undrar då hur allvarlig mintillstånd är. Detta recept är märkt `ingen påfyllnad '".
		-- Dave Barry, "Stay Fit & Healthy Until You're Dead"

%
En läkare kallar sin patient för att ge honom resultaten av hans tester. "Jag harnågra dåliga nyheter ", säger doktorn," och några sämre nyheter. "Den dåliga nyheten äratt du bara har sex veckor kvar att leva. ""Åh, nej", säger patienten. "Vad skulle kunna vara värre än det?""Jo", läkaren svarar: "Jag har försökt att nå dig sedani måndags."
		-- Dave Barry, "Stay Fit & Healthy Until You're Dead"

%
En kvinna läkare har gjort ett uttalande att rökning är varkenfysiskt defekt eller moraliskt förnedrande, och att nikotin, ävennär bortskämd i överskott, är mindre skadligt än överdriven petting. "
		-- Purdue Exponent, Jan 16, 1925

%
En kvinna gick in i ett sjukhus en dag för att föda. Efteråt läkarenkom till henne och sade: "Jag har en del ... udda nyheter för dig.""Är mitt barn okej?" frågade kvinnan oroligt."Ja, han är" doktorn svarade: "men vi vet inte hur. Din son(Vi antar) föddes med ingen kropp. Han har bara ett huvud. "Jo, doktorn var korrekt. Chefen var levande och väl, men ingenvisste hur. Chefen visade sig vara ganska normal, ignorerar hans brist påen kropp, och levde under en tid som typiskt liv som kunde förväntas enligtomständigheterna.En dag, ungefär tjugo år efter den ödesdigra födelse, kvinnan fick entelefonsamtal från en annan läkare. Läkaren sa, "Jag har nyligen fulländaten operation. Din son kan leva ett normalt liv nu: vi kan ympa en kropp påhans huvud!"Kvinnan, praktiskt gråt med glädje tackade läkaren och hängdeupp. Hon sprang uppför trappan säger, "Johnny, Johnny, har jag en * underbart *överraskning för dig! ""Åh nej," ropade Chefen, "inte en annan hatt!"
		-- Purdue Exponent, Jan 16, 1925

%
Efter hans ben hade brutits i en olycka, Mr Miller stämd för skador,claming att han var förlamad och skulle behöva tillbringa resten av sitt livi en rullstol. Även om försäkringsföretaget läkare vittnade om att hansben hade läkt ordentligt och att han var fullt kapabel att promenader,Domaren beslutade för käranden och gav honom $ 500.000.När han rullades in försäkringskassan att samla sin kontroll,Miller konfronterades av flera chefer. "Du får inte bort meddetta Miller ", en sa." Vi kommer att titta på dig dag och natt. om duta ett enda steg, kommer du inte bara återbetala skador men inför rätta förmened. Här är pengarna. Vad tänker ni göra med det? ""Min fru och jag kommer att resa", svarade Miller. "Vi ska gå tillStockholm, Berlin, Rom, Aten och slutligen till en plats som heter Lourdes -där, mina herrar, ser du er en fan av ett mirakel. "
		-- Purdue Exponent, Jan 16, 1925

%
Efter tolv års behandling min psykiater sa något somförde tårar till mina ögon. Han sa: "Nej hablo Inglés."
		-- Ronnie Shakes

%
Den som går till en psykiater borde ha huvudet undersökt.
		-- Samuel Goldwyn

%
Akvavit anses också vara användbar för medicinska ändamål, en viktigingrediens i vad jag en gång berättade är den norska botemedel för den gemensammakall. Du får en flaska, en himmelssäng, och den ljusaste färgade strumpancap du kan hitta. Du sätter locket på stolpen vid foten av sängen,sedan komma in i sängen och dricka brännvin tills du inte kan se locket. jag haraldrig provat detta, men det låter som om det borde fungera.
		-- Peter Nelson

%
Som en tumregel, aldrig lita på någon som har varit i terapiför mer än 15 procent av sin livslängd. Orden "Jag är ledsen" och "Iär fel "kommer att ha helt försvunnit från sitt ordförråd. De kommer att stickadig, skjuta dig, ha sönder saker i lägenheten, säger hemska saker till dinvänner och familj, och sedan motivera denna motbjudande beteende genom att säga:"Visst, jag sätter din hund i mikrovågsugn. Men jag känner * bättre * för att göra det."
		-- Bruce Feirstein, "Nice Guys Sleep Alone"

%
På sjukhuset, är en läkare att utbilda en praktikant på hur att meddela dåliga nyhetertill patienterna. Läkaren berättar intern "Den här mannen i 305 kommer attdö i sex månader. Gå in och tala om för honom. "Praktikanten går djärvt in irum, över till mannens BEDISDE och säger till honom "Verkar som om du kommer att dö!"Mannen har en hjärtattack och rusade in på operation på plats. DoktornGriper praktikanten och skriker på honom, "Vad!?!? är du en slags idiot?Du har att ta det lugnt, arbeta dig upp till ämnet. Nu den här mannen i213 har ungefär en vecka att leva. Gå in och tala om för honom, men försiktigt, hör du mig,försiktigt!"Praktikanten går mjukt in i rummet, humming för sig själv, cheerilyöppnar draperier att låta solen i, går över till mannens säng, luddkudden och önskar honom en "God morgon!" "Underbar dag, något att säga ...?gissa vem som kommer att dö snart! "
		-- Bruce Feirstein, "Nice Guys Sleep Alone"

%
Vara en bättre psykiater och världen kommer att slå en psykopat till din dörr.
		-- Bruce Feirstein, "Nice Guys Sleep Alone"

%
Bättre att använda läkemedel i början än i sista stund.
		-- Bruce Feirstein, "Nice Guys Sleep Alone"

%
Vissa gamla män föredrar att stiga i gryningen, med ett kallt bad och en långgå med en tom mage och i övrigt mortifying köttet. Depeka med stolthet att dessa metoder som orsaken till deras robustahälsa och mogna år; sanningen är att de är rikliga och gamla,inte på grund av sina vanor, men trots dem. Anledningen till att vi finnerbara robusta personer som utför denna sak är att det har dödat allaandra som har provat det.
		-- Ambrose Bierce, "The Devil's Dictionary"

%
Bota sjukdomen och döda patienten.
		-- Francis Bacon

%
Döden har visat sig vara 99% dödlig i laboratorieråttor.
		-- Francis Bacon

%
Tandhälsa är bredvid psykisk hälsa.
		-- Francis Bacon

%
Någonsin märker att ordet "terapeut" bryts ned till "våldtäktsmannen"?Enkel tillfällighet?Kanske...
		-- Francis Bacon

%
För min son, Robert, är detta visar sig vara hög punkten för hela sitt livhittills. Han har haft sin pyjamas på för två, kanske tre dagar nu. Han harkänslan av glädje oberoende 5-åriga barn får när han plötsligtinser att han kan driva en acetylen fackla i pälsen garderobenoch ingen av föräldrarna [på grund av influensa] skulle ha styrkan att invända.Han har födosök för sin egen mat, vilket innebär att hans diet bestårhelt av "mat" ämnen som annonseras endast på lördag morgonentecknad visar; ämnen som är färgen på jukebox ljus och att, förjuridiska skäl har deras namn felstavat, som i New CreemyChok-'n'-Cheez klumpar o 'Froot ( "en del av denna fullständiga frukost").
		-- Dave Barry, "Molecular Homicide"

%
Fortunes Motion sanningar:1: Richard Simmons får betalt för att utöva som en galning. Du behöver inte.2. Aerobic övningar stimulera och påskynda hjärtat. Så gör hjärtinfarkt.3. Träning runt små barn kan ärr dem känslomässigt för livet.4. svettas som en gris och kippar efter andan är inte uppfriskande.5. Oavsett vad någon säger, isometriska övningar kan inte göras    tyst vid skrivbordet på jobbet. Folk kommer att misstänka maniska tendenser som    du twitter runt i din stol.6. Bredvid begrava ben, saken en hund har mosts snubblar joggare.7. Låsning fyra personer i en liten, cement väggar rum så att de kan springa runt    för en timme krossa en liten gummikula - och varandra - med en hård    racket bör omedelbart erkännas för vad det är: en form av vansinne.8. Femtio armhävningar, följt av trettio sit-ups, följt av tio chin-ups,    följt av ett kast-up.9. All verksamhet som inte kan göras medan rökning bör undvikas.
		-- Dave Barry, "Molecular Homicide"

%
[Ur ett tillkännagivande av en kongress International OntopsychologyFöreningen i Rom]:Den Ontopsychological skola, som begagnar sig av nya forskningskriterier ochav en ny telematik epistemologi hävdar att sociala lägen inte vårenfrån dialektik territorium eller av klass, eller av konsumentvaror, eller medelmakt, utan snarare från dynamiska latenser capillarized i miljonerindivider i systemfunktioner som, när de väl har nått den händelsemognad, brast ut i katastrofala fenomenologi ingrepp med en lämpligstereotyp huvudpersonen eller tull marionett (allmänt, president, politiskparti, etc.) för att fullborda den handling av social schizofreni i folkmord.
		-- Dave Barry, "Molecular Homicide"

%
Gud är död och jag känner mig inte alltför väl antingen ....
		-- Ralph Moonen

%
"God hälsa" är endast den långsammaste hastigheten med vilken en kan dö.
		-- Ralph Moonen

%
Lycka är god hälsa och dåligt minne.
		-- Ingrid Bergman

%
Hälsa är bara den lägsta möjliga hastigheten med vilken man kan dö.
		-- Ingrid Bergman

%
Hälso nötter kommer att känna sig dum dag, liggande på sjukhus dörav ingenting.
		-- Redd Foxx

%
Hans idéer om första hjälpen gått så långt som sprutar sodavatten.
		-- P. G. Wodehouse

%
Humant hjärtkateterisering infördes av Werner Forssman 1929.Ignorera hans chef avdelning, och binda hans assistent en rörelsetabell för att hindra henne störningar, placerade han en uretär kateter ien ven i armen, avancerade till höger förmak [hans hjärta], ochgick uppför trapporna till röntgenavdelning där han tog bekräftanderöntgenfilm. 1956, Dr. Forssman Nobelpriset.
		-- P. G. Wodehouse

%
Jag får min motion egenskap pallbearer till mina vänner som tränar.
		-- Chauncey Depew

%
Jag fick betala för min operation. Nu vet jag vad dessa läkare varmasker för.
		-- James Boren

%
"Jag håller ser fläckar framför mina ögon.""Har du någonsin se en läkare?""Nej, fläckar bara."
		-- James Boren

%
Om en person (a) är dåligt, (b) får behandling syftar till att göra honom bättre,och (c) blir bättre, då ingen kraft resonemang känt att den medicinska vetenskapen kanövertyga honom om att det inte kan ha varit den behandling som återställde hans hälsa.
		-- Sir Peter Medawar, "The Art of the Soluble"

%
Om jag kyssa dig, är det en psykologisk interaktion.Å andra sidan, om jag slår dig i huvudet med en tegelsten,som också är en psykologisk interaktion.Skillnaden är att man är vänlig och den andra är inteså vänligt.Den springande punkten är om du kan tala om vilken som är vilken.
		-- Dolph Sharp, "I'm O.K., You're Not So Hot"

%
Om du ser ut som din körkort foto - se en läkare.Om du ser ut som din passfoto - det är för sent för en läkare.
		-- Dolph Sharp, "I'm O.K., You're Not So Hot"

%
Det är mycket vulgärt att prata som en tandläkare när en inte är en tandläkare.Det ger ett falskt intryck.
		-- Oscar Wilde.

%
Det är inte längre en fråga om att hålla sig frisk. Det är en fråga om att hittaen sjukdom som du vill.
		-- Jackie Mason

%
Det är inte verkligheten eller hur du uppfattar saker som är viktigt - det ärvad du tar för det ...
		-- Jackie Mason

%
Bara för att din läkare har ett namn för ditt tillstånd betyder inte hanvet vad det är.
		-- Jackie Mason

%
Laetrile är gropar.
		-- Jackie Mason

%
Min doktorsexamen är i litteratur, men det verkar vara en ganska bra puls till mig.
		-- Jackie Mason

%
Neurotiker bygga slott i himlen,Psykotiska lever i dem,Och psykiatriker samla hyran.
		-- Jackie Mason

%
Aldrig gå till en läkare vars kontor växter har dött.
		-- Erma Bombeck

%
New England liv, naturligtvis. Varför frågar du?
		-- Erma Bombeck

%
sida 46... En rapport citerar en studie av Dr Thomas C. Chalmers, av Mount SinaiMedical Center i New York, som jämförde två grupper som användsatt testa teorin att askorbinsyra är en kall förebyggande. "Gruppenpå placebo som trodde att de var på askorbinsyra ", säger Dr Chalmers,"Hade färre förkylningar än gruppen på askorbinsyra som trodde att de varpå placebo. "sida 56Placebo är ett bevis på att det inte finns någon verklig åtskillnad mellan kropp och själ.Sjukdom är alltid ett samspel mellan båda. Det kan börja i sinnet ochpåverka kroppen, eller den kan börja i kroppen och påverkar sinnet, som bådasom betjänas av samma blodomloppet. Försök att behandla de flesta mentalasjukdomar som om de var helt fria från fysiska orsaker och försökatt behandla de flesta kroppsliga sjukdomar som om sinnet var på något sätt inblandade måsteanses arkaiska i ljuset av nya bevis om hur människankroppsfunktioner."Anatomi av en sjukdom som uppfattas av patienten"
		-- Norman Cousins,

%
Förlamning genom analys.
		-- Norman Cousins,

%
Rätt behandling kan bota en förkylning i sju dagar, men lämnade till sig själv,en kall kommer att hänga på en vecka.
		-- Darrell Huff

%
Psykiatrin kan vi korrigera våra fel genom att bekänna våra föräldrar "brister.
		-- Laurence J. Peter, "Peter's Principles"

%
Psyko är att psykisk sjukdom som den ser sig själv en behandling.
		-- Karl Kraus

%
Psykiatri är att ta hand om id av udda.
		-- Karl Kraus

%
Visa mig en frisk människa och jag kommer att bota honom för dig.
		-- C. G. Jung

%
Psykologi. Mind over materien. Sinne i fråga? Det spelar ingen roll.Det är ingen fara.
		-- C. G. Jung

%
Pushing 30 är utöva tillräckligt.
		-- C. G. Jung

%
Pushing 40 är utöva tillräckligt.
		-- C. G. Jung

%
Sluta oroa dig för din hälsa. Det kommer att försvinna.
		-- Robert Orben

%
Sigmund hustru bar freudiansk felsägning.
		-- Robert Orben

%
Vissa människor behöver en bra imaginär botemedel mot sin smärt imaginär sjukdom.
		-- Robert Orben

%
Ibland är det bästa medicinen är att sluta ta något.
		-- Robert Orben

%
Halm? Nej, för dum en modefluga. Jag satte sot på vårtor.
		-- Robert Orben

%
Stress har lyfts fram som en viktig orsak till sjukdom. För att undvika överbelastningoch utbrändhet, hålla stressen i ditt liv. Ge den till andra i stället. Lära sigden "Gasljus" behandling, "Pratar du med mig?" teknik, och"Känner du dig okej? Du ser blek." närma sig. Börja med förhandling ochinblandning. Advance till manipulation och förnedring. Framför allt, slappna avoch ha en trevlig dag.
		-- Robert Orben

%
80-talet - när du inte kan berätta frisyrer från kemoterapi.
		-- Robert Orben

%
"... Mayo Clinic, uppkallad efter sin grundare, Dr. Ted Clinic ..."
		-- Dave Barry

%
"Kindtänderna, jag är säker på kommer att bli bra, kan molarer ta hand omsjälva ", sa den gamle mannen inte längre för mig." Men vad kommer att bliav de bicuspids? "
		-- The Old Man and his Bridge

%
New England Journal of Medicine rapporterar att nio av tio läkare är överensatt en av tio läkare är en idiot.
		-- The Old Man and his Bridge

%
Det verkliga skälet psykologi är svårt är att psykologer försökergöra det omöjliga.
		-- The Old Man and his Bridge

%
Anledningen till att de är kallade visdomständerna är att erfarenheten gör dig klok.
		-- The Old Man and his Bridge

%
Hemligheten med friska hitchhiking är att äta skräpmat.
		-- The Old Man and his Bridge

%
Problemet med hjärtsjukdom är att det första symptomet är ofta svårt attta itu med: död.
		-- Michael Phelps

%
Vet Vem Förvånad en koUnder sina uppgifter i augusti 1977 en holländsk veterinärkirurg krävdes för att behandla en sjuk ko. För att undersöka dess inregaser han införas en slang i den änden av djuret inte i stånd att ansiktsuttryck och slog en match. Strålen av eld satte eld först i visshöbalar och sedan till hela gården orsaka skador uppskattning på L45,000.Veterinären senare böter L140 för att starta en brand på ett sätt som överraskande attmagistrat. Kon undan med chock.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Vi har influensa. Jag vet inte om denna stam har en officiellnamn, men om det gör det, måste det vara något i stil med "Martian Death Flu". Dukan ha haft det själv. Det vanligaste symtomet är att du önskar att du hade en annaninställning på din elektrisk filt, upp förbi "HIGH", som sa "ELEKTRISK".Ett annat symptom är att du slutar borsta tänderna, eftersom (a)tänderna ont, och (b) du saknar styrka. Halvvägs genom borstprocess, skulle du behöva ligga ner i sink att vila ett partimmar, skulle och rännilar av tandkräm skum dribbla sidled av dinmun, så småningom härdning i knaprig lite tandkräm stalagmiter somskulle binda huvudet permanent till golvet badrum, som är hurpolisen skulle hitta dig.Du vet vilken typ av influensa jag talar om.
		-- Dave Barry, "Molecular Homicide"

%
"Välkommen tillbaka till dig 13th veckan i följd, Evelyn. Evelyn kommerdu går in i självsuggestion monter och ta din vanliga plats påpsyko-prompter soffa? ""Tack, Red.""Nu, Evelyn, förra veckan du gick upp till $ 40.000 genom att korrekt citeradin rivalitet med syskon som en tvångsmässig sado-masochistiska beteendemönster som utvecklats ur en tidig postnatal matningsproblem. ""Ja, Red.""Men - senare, när frågan om pre-adolescent oidipala fantasiförtryck, rationaliseras du två gånger och mentala blockerade tre gånger. Nu,på $ 300 per rationalisering och $ 500 per mental blocket du förlorat $ 2100 offdin $ 40,000 vilket ger ett totalt $ 37.900. Nu, någon kombination avytterligare två mentala blockeringar och antingen en rationalisering eller tre defensivaprognoser kommer att sätta dig ur spelet. Är du villig att gå vidare? ""Ja, Red.""Jag kan säga här att alla Evelyn frågor och svar harkontrollerats för noggrannhet med sin analytiker. Nu, Evelyn, för $ 80.000förklara misslyckandet med dina tre äktenskap. ""Jo, Jag--""Vi återkommer till Evelyn i en minut. Först ett ord om vårprodukt."
		-- Jules Feiffer

%
När en hel del åtgärder föreslås för en sjukdom, innebär att det inte kanbotas.
		-- Anton Chekhov, "The Cherry Orchard"

%
Matsmältningssystemet är kroppens Fun House, där mat går på en lång,mörk, skrämmande rida, ta alla typer av oväntade vändningar, ärattackeras av onda sekret längs vägen, och inte veta till sistaminut om det kommer att förvandlas till en användbar kroppsdel ​​eller sprutas in iMörkt hål av Mister Sfinkter. Vi amerikaner lever i en nation därmedicinsk-och sjukvårdssystemet är oöverträffad i världen, om man räknar kanske25 eller 30 små scuzzball länder som Skottland som vi kunde förångas isekunder om vi kändes som det.
		-- Dave Barry, "Stay Fit & Healthy Until You're Dead"

%
