Steg 1: Stäng AutoCAD - Jag vet att det kan vara svårt för vissa av er. Du kundeockså vänta för AutoCAD att krascha om du vill.    - Michael Rotolo       (Http://themadcadder.blogs.com/my_weblog/2008/12/external-xref-manager-xref-path-saver.html)! 11/07 PDP en Ni deppart m'I! PleH
		-- Jamie Zawinski

%
101 ANVÄNDNING SFOR En död MIKROPROCESSOR(1) Scarecrow för tusenfotingar(2) Dead katt borste(3) Hår barrettes(4) Inre stöd(5) Själv piercing örhängen(6) Fungus spaljé(7) Lösögonfransar(8) Prosthetic hund klorna        .        .        .(99) Fönster trädgård harv (dras bakom Tonka traktorer)(100) Killer velcro(101) Valuta
		-- Jamie Zawinski

%
1: Ingen kodtabell för OP: ++ post
		-- Jamie Zawinski

%
4,2 BSD UNIX # 57: Sun 1 juni 23:02:07 EDT 1986Du svänga på solen Du saknar. Solen svänger. Han slår dig med en575MB disk! Du läser 575MB disk. Den är skriven på ett främmandetunga och kan inte läsas av dina trötta Sun-2 ögon. Du kastar575MB skivan vid sön Du träffar! Solen måste reparera dina ögon. DeSun läser en scroll. Han slår din 130 MB disk! Han har besegrat130 MB disk! Solen läser en scroll. Han träffar din Ethernet-kortet! hanhar besegrat din Ethernet-kortet! Du läser en rulla av "skjuta framMåndag klockan 09:00 ". Allting går mörkt ...
		-- /etc/motd, cbosgd

%
En biolog, en statistiker, en matematiker och datavetare är påen fotosafari i Afrika. När de kör längs savannen i derasjeep, de stannar och spana horisonten med sina kikare.Biologen: "Titta En flock av zebror Och det finns en vit zebra!!	Fantastisk! Vi ska vara känd! "Statistikern: "Hej, lugna ner, det är inte signifikant Vi vet bara.Det finns en vit zebra. "Matematikern: "Egentligen är vi bara vet att det existerar en zebra, som ärvit på ena sidan. "Datorn forskare: "Åh nej Ett specialfall!"
		-- /etc/motd, cbosgd

%
... En blomstrande röst säger: "Fel, cretin!", Och du märker att duhar förvandlats till en hög av damm.
		-- /etc/motd, cbosgd

%
Ett fel i koden är värt två i dokumentationen.
		-- /etc/motd, cbosgd

%
Ett fel i handen är bättre än en ännu oupptäckt.
		-- /etc/motd, cbosgd

%
En viss munk hade en vana av tjat Grand Tortue (den enda somnågonsin nått upplysningen "Yond upplysningen), genom att fråga omolika objekt hade Buddha-natur eller inte. På en sådan fråga Tortuealltid satt tyst. Munken hade redan bett om en böna, en sjö,och en månbelyst natt. En dag han förde till Tortue ett snöre, ochställde samma fråga. Som svar, Grand Tortue fattade slinganmellan hans fötter och, med några få enkla handgrepp, skapade en komplexsträng som han proferred wordlessly till munken. I det ögonblicket, munkenvar upplyst.Från och med då, gjorde munken inte bry Tortue. Istället gjorde han sträng eftersträngen genom Tortue metod; och han passerade metoden vidare till sina egna elever,som passerade den på till deras.
		-- /etc/motd, cbosgd

%
Ett komplext system som fungerar är alltid visade sig ha utvecklats från enenkelt system som fungerar.
		-- /etc/motd, cbosgd

%
[En dator är] som en gammaltestamentlig gud, med en mängd regler och ingen nåd.
		-- Joseph Campbell

%
En dator kan du göra fler misstag snabbare än någon annan uppfinning,med eventuella undantag för handeldvapen och Tequilla.
		-- Mitch Ratcliffe

%
En dator försäljare besöker en vd för att säljaordföranden en av de senaste talande datorer.Säljare: "Den här maskinen vet allt jag kan ställa det någon fråga.och det kommer att ge det rätta svaret. Dator, vad är		ljusets hastighet?"Dator: 186,282 miles per sekund.Säljare: "Vem var den första presidenten i USA?"Dator: George Washington.Ordförande: "Jag är fortfarande inte övertygad Låt mig ställa en fråga..Var är min far? "Dator: Din far fiskar i Georgien.Ordförande: "Hah !! Datorn är fel Min far dog över tjugo.		för flera år sedan!"Dator: Din mor make dog för 22 år sedan. Din far baralandade en tolv pund bas.
		-- Mitch Ratcliffe

%
En datavetare är någon som fixar saker som inte är trasiga.
		-- Mitch Ratcliffe

%
En dator utan COBOL och Fortran är som en bit chokladkakautan ketchup och senap.
		-- Mitch Ratcliffe

%
En CONS är ett föremål som bryr sig.
		-- Bernie Greenberg.

%
Ett debuggade program är ett som du ännu inte har hittat de villkorsom gör det misslyckas.
		-- Jerry Ogdin

%
En lärjunge till en annan sekt gång kom till Drescher som han äterhans morgonen måltid. "Jag skulle vilja ge dig den här personlighetstest", sadeutomstående ", eftersom jag vill att du ska vara lycklig."Drescher tog det papper som erbjöds honom och placera den ibrödrost - "Jag önskar brödrosten att vara glad för."
		-- Jerry Ogdin

%
En läkare, en arkitekt, och datavetare grälade omvars yrke var den äldsta. Under sina argument, defick hela vägen tillbaka till Edens lustgård, varpå läkaren sa, "läkarkåren är klart den äldsta, eftersom Eva gjordes från Adamsrevben, som historien går, och det var en helt enkelt otroligt kirurgisk bedrift. "Arkitekten inte överens. Han sa: "Men om man tittar på Gardensjälv, i början var det kaos och ogiltiga, och ur den trädgårdenoch världen skapades. Så Gud måste ha varit en arkitekt. "Den datorforskare, som hade lyssnat noga på allt detta, dåkommenterade: "Ja, men där tror ni kaoset kom ifrån?"
		-- Jerry Ogdin

%
En känd Lisp Hacker märkte en Grundutbildning sitter framför en Xerox1108, försöker redigera ett komplext Klone nätverk via en webbläsare. viljahjälp, Hacker klickade en av noderna i nätverket med musen,och frågade "Vad ser du?" Mycket allvarligt, svarade Grundutbildning "Jagse en markör. "The Hacker sedan snabbt tryckte på start växla på baksidanpå tangentbordet och samtidigt trycka på Undergraduate över huvudetmed en tjock Interlisp Manual. Student var sedan upplyst.
		-- Jerry Ogdin

%
En formell tolkning algoritm inte alltid användas.
		-- D. Gries

%
En Fortran kompilator är troll av små minis.
		-- D. Gries

%
En hacker gör för kärlek vad andra inte skulle göra för pengarna.
		-- D. Gries

%
Ett språk som inte påverkar ditt sätt att tänka om programmering ärinte värt att veta.
		-- D. Gries

%
Ett språk som inte har allt är faktiskt lättare att programmerai än vissa som gör det.
		-- Dennis M. Ritchie

%
Ett stort antal installerade system fungerar genom fiat. Det vill säga, de arbetargenom att ha deklarerats arbeta.
		-- Anatol Holt

%
En LISP programmerare vet värdet av allt, men kostnaden för ingenting.
		-- Alan Perlis

%
En lista är inte starkare än sin svagaste länk.
		-- Don Knuth

%
En liten tillbakablickande visar att även om många fina, användbara mjukvarusystemhar utformats av utskotten och byggdes som en del av flera delar projekt,dessa mjukvarusystem som har glada passionerade fans är de som ärprodukter från en eller ett fåtal utforma sinnen, stora designers. Överväga Unix,APL, Pascal, Modula, Smalltalk-gränssnittet, även Fortran; och kontras demmed Cobol, PL / I, Algol, MVS / 370, och MS-DOS.
		-- Fred Brooks

%
En man från AI gick över bergen för att segla till se Master,Knuth. När han kom, Mästaren var ingenstans att hittas. "Var ärklokt som heter Knuth? "frågade han en förbipasserande student."Ah", sade studenten, "du inte har hört. Han har gått på enpilgrimsfärd över bergen till templet i AI att söka nyalärjungar. "Hörde detta, var mannen upplyst.
		-- Fred Brooks

%
En chef frågade en programmerare hur lång tid det skulle ta honom att avslutaprogram som han arbetade. "Jag kommer att vara klar i morgon," programmerarenomgående svarade."Jag tror att du är orealistiska", sade chefen. "Sanningsenligt,hur lång tid tar det?"Programmeraren trodde för ett ögonblick. "Jag har några funktioner som jag villtillägga. Detta kommer att ta minst två veckor, "äntligen sade han."Även det är för mycket att förvänta sig", insisterade chefen, "Jag kommer att varanöjd om du helt enkelt tala om för mig när programmet är klart. "Programmeraren gick med på detta.Flera år senare, pensionerad chef. På väg till sinpension lunch upptäckte han programmeraren sover vid sin terminal.Han hade programmering hela natten.
		-- Geoffrey James, "The Tao of Programming"

%
En chef var på väg att få sparken, men en programmerare som arbetade för honomuppfann ett nytt program som blev populär och sålde bra. Som ett resultat, denmanager behöll sitt jobb.Chefen försökt att ge programmeraren en bonus, men programmerarenvägrade det, säger, "jag skrev programmet eftersom jag att det var en intressantkoncept, och därför förväntar jag mig ingen belöning. "Chefen, när han hörde detta, sade: "Detta programmerare, men hanhar en ställning av små känsla, förstår väl rätt plikt enanställd. Låter befordra honom till upphöjd position managementkonsult! "Men då berättade detta, programmeraren gång vägrade och sade: "Jag existerarså att jag kan programmera. Om jag var främjas, skulle jag inte göra annat än avfallallas tid. Kan jag gå nu? Jag har ett program som jag arbetar på. "
		-- Geoffrey James, "The Tao of Programming"

%
En chef gick till sina programmerare och sade till dem: "När det gäller dinarbetstid: du kommer att behöva komma in på nio på morgonen och lämnavid fem på eftermiddagen. "På detta, alla av dem blev arg och fleraavgick på plats.Så chefen sade: "Okej, i så fall kan ställa in din egenarbetstid, så länge du är klar med projekt på schemat. "Detprogrammerare, nu nöjd, började komma i en middag och arbeta för att pissamorgontimmarna.
		-- Geoffrey James, "The Tao of Programming"

%
En chef gick till huvudprogrammerare och visade honom de kravdokumentera för en ny ansökan. Chefen frågade befälhavaren: "Hur länge kommerdet tar att utforma detta system om jag tilldelar fem programmerare till det? ""Det kommer att ta ett år", sade befälhavaren omgående."Men vi behöver detta system omedelbart eller ens förr! Hur lång tid tar detta det tilldelar jag tio programmerare till det? "Befälhavaren programmerare rynkade pannan. "I så fall kommer det att ta två år.""Och om jag tilldela hundra programmerare till det?"Befälhavaren programmerare lättvindigt. "Då designen kommer aldrig att blifärdig ", sade han.
		-- Geoffrey James, "The Tao of Programming"

%
En mästare programmerare passerade en novis programmerare en dag. Mästarennoterade nybörjare upptagenhet med en handhållen dataspel. "Ursäkta mig",sade han, "kan jag undersöka det?"Novisen bultad till uppmärksamhet och överlämnade enheten till master."Jag ser att enheten påstår sig ha tre nivåer av spel: Lätt, Medium,och hårt ", sade befälhavaren." Men varje sådan anordning har en annan nivå av lek,där anordningen försöker inte att erövra människors eller att besegras avmänsklig.""Be, store mästare" bad novisen, "hur man hittarmystisk inställning? "Befälhavaren tappade enheten till marken och krossade den under fötterna.Och plötsligt nybörjare var upplyst.
		-- Geoffrey James, "The Tao of Programming"

%
En master förklarade natur Tao till ett av sina nybörjare."Tao förkroppsligas i alla program - oavsett hur obetydlig"sade befälhavaren."Är Tao i en handhållen miniräknare?" frågade nybörjare."Det är" kom svaret."Är Tao i ett videospel?" fortsatte nybörjare."Det är ännu i ett videospel," sade befälhavaren."Och är Tao i DOS för en personlig dator?"Befälhavaren hostade och skiftade sin position något. "Lektionenär över för i dag ", sade han.
		-- Geoffrey James, "The Tao of Programming"

%
Ett modem är en Baudy hus.
		-- Geoffrey James, "The Tao of Programming"

%
En otäck snygga dvärg kastar en kniv på dig.
		-- Geoffrey James, "The Tao of Programming"

%
*** En ny typ av programmering ***Vill du omedelbar respekt som kommer från att kunna använda teknisktermer som ingen förstår? Vill du sätta skräck och avsky ihjärtan DP chefer överallt? Om så är fallet, låt den berömda programmerare "Skola leda dig på ... i en värld av professionell datorprogrammering.De säger att en bra programmerare kan skriva 20 rader effektivt program per dag.Med vår unika utbildning, så visar vi dig hur man skriver 20 rader kodoch mycket annat. Vår utbildning täcker alla programmeringsspråkexisterar, och några som inte är det. Du lär dig varför on / off knapp för endator är så viktigt, vad orden * allvarligt fel * betyder, och vem och vaddu bör skylla på när du gör ett misstag.Ja, jag vill broschyr som beskriver denna otroliga erbjudande.Jag bifogar $ 1000 är små omärkta räkningar för att täcka kostnaderna förporto och hantering. (Inga levande fjäderfän, tack.)*** Vår slogan: Top down programmering för massorna. ***
		-- Geoffrey James, "The Tao of Programming"

%
En novis frågade Mästaren: "Här är en programmerare som aldrig designar,dokument, eller tester hans program. Men alla som känner honom betraktar honom en avde bästa programmerare i världen. Varför är detta?"Mästaren svarar: "Det programmerare har bemästrat Tao Han har.gått utöver behovet av design; Han blir inte arg när systemetkraschar, men accepterar universum utan bekymmer. Han har gått längre änbehovet av dokumentation; han inte längre bryr sig om någon annan ser sin kod. hanhar gått längre än nödvändigt för att testa; vart och ett av hans program är perfekt inomsjälva, lugn och elegant, deras syfte självklart. Sannerligen, har hanin i mysteriet med Tao. "
		-- Geoffrey James, "The Tao of Programming"

%
En novis frågade befälhavaren: "Jag har ett program som ibland körs ochibland avbryts. Jag har följt reglerna för programmering, men jag är heltsnopen. Vad är orsaken till detta? "Befälhavaren svarade: "Du är förvirrad eftersom du inte förstårTao. Bara en dåre förväntar rationellt beteende från sina medmänniskor. Varförförväntar du dig det från en maskin som människor har konstruerat? datorersimulera determinism; bara Tao är perfekt.Reglerna för programmering är övergående; bara Tao är evig.Därför måste du överväga Tao innan du får upplysning. ""Men hur vet jag när jag har fått upplysning?" frågadenybörjare."Ditt program kommer då att fungera", svarade befälhavaren.
		-- Geoffrey James, "The Tao of Programming"

%
En novis frågade befälhavaren: "Jag upplever att ett dataföretag ärmycket större än alla andra. Det höjer sig över dess konkurrens som en gigantiskbland dvärgar. Vilken som helst av dess divisioner kan innefatta en hel verksamhet.Varför är det så? "Befälhavaren svarade: "Varför frågar du så dumma frågor? Detföretag är stor eftersom det är så stor. Om det bara gjort hårdvara, ingenskulle köpa den. Om det bara underhållna system, skulle människor behandlar det som entjänare. Men eftersom den kombinerar alla dessa saker, människor tycker att det enav gudarna! Genom att inte försöka sträva, erövrar det utan ansträngning. "
		-- Geoffrey James, "The Tao of Programming"

%
En novis frågade befälhavaren: "I öster finns en stor trädstrukturatt män kallar "Corporate högkvarter". Det är uppsvälld ur form medvice ordförande och revisorer. Det ger en mängd PM, var att säga"Gå, alltså! eller "Gå, Hit! och ingen vet vad som menas. Varje år nyanamn sätts på grenarna, men alla till ingen nytta. Hur kan en sådanonaturliga enhet existerar? "Befälhavaren svarar: "Du uppfattar denna enorma struktur och ärstörd att den inte har någon rationell syfte. Kan du inte ta nöje fråndess oändliga vändningar? Tycker du inte njuta av obesvärad enkel programmeringunder dess skyddande grenar? Varför är du besväras av sin värdelöshet? "
		-- Geoffrey James, "The Tao of Programming"

%
En nybörjare i templet en gång närmade sig översteprästen med enfråga."Mästare, gör Emacs har Buddha-natur?" nybörjare frågade.Översteprästen hade varit i templet i många år och kan varaåberopas för att veta dessa saker. Han tänkte i flera minuter innansvara."Jag förstår inte varför inte. Det har fått banne allt annat."Därmed gick översteprästen till lunch. Novisen plötsligtuppnås upplysning, flera år senare.Kommentar:Hans Master är snäll,Svara hans FAQ snabbt,Med tanke och sarkasm.
		-- Geoffrey James, "The Tao of Programming"

%
En nybörjare programmerare en gång tilldelats koda en enkel finansiellpaket.Novisen arbetade ursinnigt i flera dagar, men när hans herreöver sitt program, upptäckte han att det innehöll en textredigeraren, en uppsättningAllmänna grafikrutiner och artificiell intelligens gränssnitt,men inte det minsta omnämnande av något ekonomiskt.När befälhavaren frågade om detta, blev nybörjare upprörd."Var inte så otålig", sade han, "jag ska sätta den finansiella grejer så småningom."
		-- Geoffrey James, "The Tao of Programming"

%
En nybörjare försökte fixa en trasig lisp maskinen genom att vridaströmmen och på. Knight, se vad eleven gjorde yttrade strängt,"Du kan inte fixa en maskin genom att bara power-cykling det med någon förståelseav vad som går fel. "Knight vände maskinen av och på. Denmaskin fungerade.
		-- Geoffrey James, "The Tao of Programming"

%
En person som är mer än vardag intresserad av datorer bör vara välskolad i maskinkod, eftersom det är en grundläggande del av en dator.
		-- Donald Knuth

%
Ett program bör vara lätt och smidig, dess subrutiner ansluten som ensträngar av pärlor. Andemeningen och syftet med programmet bör behållasgenom hela. Det bör varken vara för lite eller för mycket, varken onödigtslingor eller onödiga variabler, varken brist på struktur eller överväldigandestelhet.Ett program bör följa "Lagen om minst förvåning". Vad är dettalag? Det är helt enkelt att programmet alltid ska svara för användaren isätt som förvånar honom minst.Ett program, oavsett hur komplex, bör fungera som en enda enhet. DeProgrammet bör ledas av logiken i stället för genom systemet för passivutseenden.Om programmet inte i dessa krav, kommer det att vara i ett tillstånd avoordning och förvirring. Det enda sättet att rätta till detta är att skriva omprogram.
		-- Geoffrey James, "The Tao of Programming"

%
En programmerare från en mycket stor dataföretag gick till en programvarakonferens och återvände sedan rapportera till sin chef, säger: "Vad för slagsprogrammerare arbetar för andra företag? De betedde sig illa och varobekymrad med framträdanden. Deras hår var långt och misskött och deraskläder var skrynkliga och gamla. De kraschade ut gästfrihet sviter och degjort oförskämd ljud under min presentation. "Chefen sa: "Jag skulle aldrig ha skickat dig till konferensen.Dessa programmerare lever bortom den fysiska världen. De anser liv absurt,en oavsiktlig tillfällighet. De kommer och går utan att veta begränsningar.Utan en omsorg, de lever bara för sina program. Varför skulle de brymed sociala konventioner? ""De lever inom Tao."
		-- Geoffrey James, "The Tao of Programming"

%
En programmerare är en person som passerar som en krävande expert på grundval avatt kunna visa sig, efter otaliga stansning, en oändlig serie avobegripliga svar beräknade med mikrometerprecisionerna från vagaantaganden baserade på diskutabla siffror tagna från ofullständiga handlingaroch utföras på instrument problematisk noggrannhet av personer medtvivelaktiga tillförlitlighet och tveksamt mentalitet för det uttalade syftet medirriterande och blanda ihop en hopplöst försvarslös avdelning som varoturen att be om information i första hand.
		-- IEEE Grid newsmagazine

%
Ett programmeringsspråk är låg nivå när dess program kräver uppmärksamhettill irrelevant.
		-- IEEE Grid newsmagazine

%
En ny studie har funnit att koncentrera sig på svåra off-screenföremål, såsom ansikten nära och kära, orsakar påfrestningarna på ögonen i datornvetenskapsmän. Forskare i fenomenet citera den tillsatta koncentrationensom behövs för att "vettigt" av sådana onaturliga tredimensionella objekt.
		-- IEEE Grid newsmagazine

%
En rullande disk samlar ingen MOS.
		-- IEEE Grid newsmagazine

%
En student, i hopp om att förstå Lambda-karaktär, kom till Greenblatt.När de talade Multics systemet hacker promenerade genom. "Är det sant", frågadeelev "att PL-1 har många av de samma datatyper som Lisp?" nästan innaneleven hade avslutat sin fråga, Greenblatt ropade "foo", och slåstudenten med en pinne.
		-- Jack Banton, PCC Automotive Electrical School

%
En framgångsrik [programvara] verktyg är ett som användes för att göra någotoanade av dess författare.
		-- S. C. Johnson

%
En väl använt dörr behöver ingen olja på sina gångjärn.Ett snabbt strömmande ånga växer inte stillastående.Varken ljud eller tankar kan färdas genom ett vakuum.Programvaru ruttnar om den inte används.Dessa är stora mysterier.
		-- Geoffrey James, "The Tao of Programming"

%
Ett år tillbringade i artificiell intelligens är tillräckligt för att få en tro på Gud.
		-- Geoffrey James, "The Tao of Programming"

%
Om användningen av språket: det är omöjligt att vässa en penna med en trubbigyxa. Det är lika fåfängt att försöka göra det med tio trubbiga axlar i stället.
		-- Edsger Dijkstra

%
Lägga till funktioner inte nödvändigtvis öka funktionaliteten - det baragör handböckerna tjockare.
		-- Edsger Dijkstra

%
Lägga arbetskraft till en sen programvaruprojekt gör det senare.
		-- F. Brooks, "The Mythical Man-Month"

%
När en person befinns lämpligt för utsläpp av en skyldighet avStäng programmet därtill, är det värre köra med två personer ochknappast gjort alls om tre eller fler anställda däri.
		-- George Washington, 1732-1799

%
Efter siktning genom de skrivna återstående block av Luke hemkatalog, Luke och PDP-1 accelererade bort från / u / Lars, över ytan på denWinchester ridning Lukes flygande läs / skrivhuvudet. PDP-1 hade Luke stopp vidkanten av cylindern med utsikt / usr / spool / uucp."Unix-till-Unix Copy Program;" sade PDP-1. "Du kommer aldrig hitta en merusel sjuder av buggar och flamers. Vi måste vara försiktiga. "
		-- DECWARS

%
Alan Turing tänkte om kriterier för att lösa frågan ommaskiner kan tänka, en fråga som vi nu vet att det handlar omså relevant som frågan om ubåtar kan simma.
		-- Dijkstra

%
Algol-60 säkert måste betraktas som den viktigaste programmeringsspråkännu inte utvecklat.
		-- T. Cheatham

%
Alla konstanter är variabler.
		-- T. Cheatham

%
=== ALLA CSH ANVÄNDARE OBS ========================Ställ in variabeln $ FÖRLORARE till alla de människor som du tycker är förlorare. Dettakommer att orsaka alla dessa förlorare har variabeln $ PEOPLE-WHO-THINK-I-AM-A-FÖRLORAREuppdateras i deras .login. Om du försöker köra ett jobb på enmaskin med dålig svarstid och en maskin på din lokala nätet är för närvarandebefolkad av förlorare, kommer att maskinen frigörs för jobbet genom enkall startprocessen.
		-- T. Cheatham

%
Alla delar ska gå ihop utan att tvinga. Du måste komma ihåg att de delardu återmontering var demonteras av dig. Därför, om du inte kan fåihop dem igen, måste det finnas en anledning. Med alla medel, inte använda en hammare.
		-- IBM maintenance manual, 1925

%
Alla programmerare är optimister. Kanske denna moderna trolldom särskilt lockardem som tror på ett lyckligt slut och fairy gudmödrar. Kanske hundratalsav praktiska frustration köra bort alla utom de som vanligtvis fokuserar på slutetmål. Kanske är det bara att datorer är unga, programmerare är yngre,och de unga är alltid optimister. Men hur urvalsprocessen fungerarResultatet är odiskutabelt: "Den här gången kommer säkert köra" eller "Jag hittadeden sista felet. "
		-- Frederick Brooks, "The Mythical Man Month"

%
Alla programmerare är dramatiker och alla datorer är usel skådespelare.
		-- Frederick Brooks, "The Mythical Man Month"

%
"... Alla goda data mönster bootlegged, den formellt planeradeprodukter, om de byggs alls, är hundar! "MIT Press, 1987
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
Alla de enkla program har skrivits.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================Ett nytt system, cirkulationssystemet, har lagts till.Den lång experimentella cirkulationssystemet har släppts till användarna. DeLisp Machine använder typ B vätska, använder L maskintyp En vätska. närByt till Common Lisp inträffar båda maskinerna kommer naturligtvis att vara typ O.Kontrollera vätskenivån med hjälp av oljestickan som ligger i denbaksidan av VMI monitorer. Okontrollerade låga vätskenivåer kan orsaka dålig ökningprestanda.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================Felrapporter uppgår nu till i genomsnitt 12.853 per dag. Tyvärr,Detta är bara en liten del [<1%] av postvolymen vi får. Ibesluta att vi mer skyndsamt kan ta itu med dessa värdefulla meddelandenvänligen meddela dem genom en av följande vägar:ARPA: WastebasketSLMHQ.ARPAUUCP:!!!! [Berkeley, seismo, harpo] fubar thekid slmhq papperskorg Icke-nätverksplatser: Federal Express till:papperskorgroom NE43-926Copernicus, månen, 12345-6789För att personlig kontakt känsla samtal 1-415-642-4948; vår utbildadeoperatörer har jour 24 timmar om dygnet. VISA / MC accepteras. ** Våra mycket rika jurister har försäkrat oss om att vi inte  ansvarig för eventuella fel eller råd som ges via telefon.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================BIL och CDR nu återvända extra värden.Funktionen CAR returnerar nu två värden. Eftersom det har att gå till besvärta reda på om objektet är carcdr-kan i alla fall, vi tänkte du kanske somväl få båda halvorna på en gång. Till exempel visar följande kod hur mandestrukturera en cons (något-CONS) i sina två kortplatser (THE-CAR och THE-CDR):(FLERA värde BIND (THE-bil-CDR) (CAR NÅGRA-CONS) ...)För symmetri med CAR, CDR returnerar ett andra värde som är bilen förobjekt. I en relaterad förändring, funktioner gör-array och CONS har varitfast så att de inte tilldela någon lagring utom på stacken. detta börförhoppningsvis hjälpa människor som inte gillar att använda sophämtare eftersomdet kalla stövlar maskinen så ofta.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================Kompilator optimeringar har gjorts till makro expandera LET in i en WITHOUT-INTERRUPTS speciell form så att den kan driva saker till en stapel iLET optimering området setq variablerna och sedan pop dem tillbaka när det ärgjort. Oroa dig inte om detta om du inte använder multi.Observera att LET * kunde * har definierats av:(LET ((LET '' (LET ((LET ', LET)), LET)))'(LET ((LET', LET)), LET))Detta tros påskynda utförande med så mycket som en faktor av 1,01 eller3,50 beroende på om du tror att våra vänliga marknadsföring representanter.Denna kod är skriven av en ny programmerare här (vi ryckte bort honom frånItty Bitti Machines där han skrev COUGHBOL kod) så att ge honomförtroende vi betrodda hans löften om "det fungerar ganska bra" och installerat den.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================JCL stöd som alternativ till systemmenyn.I vår fortsatta ansträngningar för att stödja andra språk än Lisp på CADDR,Vi har utvecklat ett OS / 360-kompatibel JCL. Detta kan användas som enalternativ till den vanliga systemmenyn. Typsystem J för att komma till en JCLinteraktiv skriv köra diagnostisera slingfönstret. [Notera att för 360kompatibilitet, alla ingångslinjer avkortas till 80 tecken.] Dennafönster har även en mus känslig visning av kritiska parametrar jobbsåsom dataset tilldelning, kärn tilldelning, kanaler, etc. När en JCLsyntaxfel upptäcks eller ditt jobb abends, fönsterorienterade JCLdebugger anges. Den JCL debugger visar lämplig OS / 360 felmeddelanden (såsom IEC703 "disk error") och låter dig avköa ditt jobb.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================Skräpinsamlaren fungerar nu. Dessutom en ny, experimentell soporsamling algoritm har installerats. Med SI:% DSK-GC-QLX-BITS satt till 17,(INTE standard) gamla sophämtning algoritm är i kraft; närvirtuellt minne fylls maskinen kalla stövlar själv. Med SI:% DSK-GC-QLX-bitar satta till 23, den nya sophämtare aktiverad. Till skillnad från de flesta soporsamlare, startar nya gc sin prägel fasen från minnet av användaren, snarareän från obarray. Detta gör det möjligt för sophämtning avsevärtmera Qs. Som skräpinsamlaren körs kan det fråga dig något liknande "Har duihåg vad SI: RDTBL-TRANS gör ", och om du inte kan ge ett rimligt svar?i trettio sekunder, blir symbolen en kandidat för GCing. den rörligaSI:% GC-QLX-Luser-TM styr hur länge GC väntar innan timing ut användaren.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
=== ALLA ANVÄNDARE OBS ========================Det har rått viss förvirring om MAPCAR.(Defun MAPCAR (& FUNKTIONELL FCN & EVAL och avkoppling listor)(PROG (V P LP)(Setq P (LOCF V))L (setq LP listor)(% START-FUNKTION-CALL FCN T (längd listor) NIL)L1 (OR LP (GO L2))(OCH (NULL (CAR LP)) (RETURN V))(% PUSH (caar LP))(RPLACA LP (CDAR LP))(Setq LP (CDR LP))(GO L1)L2 (% FINISH-FUNKTION-CALL FCN T (längd listor) NIL)(Setq LP (% POP))(RPLACD P (setq P (NCONS LP)))(GO L)))Vi hoppas att detta rensar upp många frågor som vi har haft om det.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
Alla dina filer har förstörts (sorry). Paul.
		-- David E. Lundstrom, "A Few Good Men From Univac",

%
Nästan allt nedsättande man kan säga om dagens mjukvarudesignskulle vara korrekt.
		-- K. E. Iverson

%
Även om det fortfarande en truism inom industrin att "ingen någonsin fick sparken förköpa IBM, "Bill O'Neil, den teknikchef på Drexel BurnhamLambert, säger att han vet för ett faktum att någon har fått sparken för just dettaanledning. Han vet det eftersom han sköt killen."Han gjorde ett dåligt beslut, och vad det kom ner till var," Ja, jagköpte det eftersom jag tänkte att det var säkert att köpa IBM, "" Mr O'Neil säger."Jag sa," Nej Fel. Game over. Nästa tävlande, tack. ""
		-- The Wall Street Journal, December 6, 1989

%
AmigaDOS Öl: Företaget har gått i konkurs, men deras recept hartagits upp av några konstiga tyska företaget, så nu detta öl kommer att vara enimportera. Detta öl aldrig riktigt sålt mycket bra eftersom den ursprungligatillverkaren inte förstår marknadsföring. Som Unix öl, AmigaDOS ölfans är en extremt lojal och högljudd grupp. Det kom ursprungligen i en16-oz. kan, men nu kommer i 32-oz. burkar också. När detta kan varursprungligen infördes, föreföll det spännande och färgstark, men designenhar inte förändrats mycket under åren, så det verkar daterad nu. kritiker avdenna öl hävdar att det endast är avsedd för att titta på TV hur som helst.
		-- The Wall Street Journal, December 6, 1989

%
Ett undantag Ada är när en rutin får problem och säger"Beam me up, Scotty".
		-- The Wall Street Journal, December 6, 1989

%
En adekvat bootstrap är en självmotsägelse.
		-- The Wall Street Journal, December 6, 1989

%
En algoritm måste ses att döma.
		-- D. E. Knuth

%
... En anekdot från IBM: s Yorktown Heights Research Center. När enprogrammerare använde sin nya datorterminal, allt var bra när han sattner, men han kunde inte logga in i systemet när han stod upp. Den därbeteende var 100 procent repeterbar: han kunde alltid logga in när man sitter ochaldrig när du står.De flesta av oss bara luta dig tillbaka och förundras över en sådan berättelse; Hur kunde det terminalvet om den stackars killen var sittande eller stående? Goda debuggers, fast,vet att det måste finnas en anledning. Elektriska teorier är lättast atthypotes: var det en lös tråd under mattan, eller problem med statiskelektricitet? Men elektriska problem är sällan genomgående reproducerbar.En varning IBMer slutligen märkte att problemet var i terminalens tangentbord:toppar två nycklar byttes. När programmeraren satt han var entouch-metoden och problemet gick obemärkt, men när han stod han leddesvilse av jakt och picka.
		-- "Programming Pearls" column, by Jon Bentley in CACM February 1985

%
En elefant är en mus med ett operativsystem.
		-- "Programming Pearls" column, by Jon Bentley in CACM February 1985

%
En ingenjör är någon som gör lista behandling i Fortran.
		-- "Programming Pearls" column, by Jon Bentley in CACM February 1985

%
En tolkning _ I uppfyller en mening i tabellen språk om och endast omvarje post i tabellen betecknar värdet av funktionen betecknad medFunktionen konstant i det övre vänstra hörnet tillämpas på objekten utseddamed motsvarande rad- och kolumnetiketter.intelligens "
		-- Genesereth & Nilsson, "Logical foundations of Artificial

%
Och det bör vara lagen: Om du använder ordet 'paradigm "utan att vetaVad ordboken säger att det betyder, du går till fängelse. Inga undantag.
		-- David Jones

%
Och på den sjunde dagen, han lämnat bifogningsläge.
		-- David Jones

%
En annan megabyte dammet.
		-- David Jones

%
Ett visst program kommer att expandera för att fylla det tillgängliga minnet.
		-- David Jones

%
Ett visst program, när du kör, är föråldrad.
		-- David Jones

%
Alla program som körs rätt är föråldrad.
		-- David Jones

%
Alla programmeringsspråk är bäst innan den genomförs och används.
		-- David Jones

%
... Alla likheter mellan ovanstående synpunkter och de min arbetsgivare,min terminal eller vyn ut mitt fönster är en ren slump. Någralikhet mellan ovanstående och mina egna åsikter är icke-deterministiska. DeFrågan om förekomsten av åsikter i avsaknad av någon att hålla demär kvar som en övning för läsaren. Frågan om det föreliggerläsaren är kvar som en övning för andra gud koefficienten. (ENdiskussion av icke-ortogonala, icke-integrerad polyteism ligger utanför rameni den här artikeln.)
		-- David Jones

%
Alla tillräckligt avancerad bugg är omöjlig att skilja från en funktion.
		-- Rich Kulawiec

%
Den som har deltagit i en USENIX konferens i ett fint hotell kan berättaatt en mening som "Du är en av dessa dator människor, eller hur?"motsvarar ungefär "Titta, en annan otroligt mobil form av slemmögel! "i munnen på ett hotell servitris.
		-- Elizabeth Zwicky

%
APL hackare gör det i quad.
		-- Elizabeth Zwicky

%
APL är ett misstag, genomföras till perfektion. Det är det språk somframtid för programmeringsteknik i det förflutna: det skapar en ny generationav kodande bums.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
APL är en naturlig förlängning av assembler programmeringsspråk;... Och är bäst för utbildningsändamål.
		-- A. Perlis

%
APL är en skriv enda språk. Jag kan skriva program i APL, men jag kan inteläst någon av dem.
		-- Roy Keir

%
Vi kör ljus med overbyte?
		-- Roy Keir

%
Runt datorer är det svårt att hitta rätt tidsenhet tillmäta framstegen. Vissa katedraler tog ett sekel att slutföra. Kan duföreställa sig storheten och omfattningen av ett program som skulle ta så lång tid?
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Som en dator, jag tycker din tro på teknik underhållande.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Såvitt vi vet har vår dator aldrig haft ett oupptäckt fel.
		-- Weisert

%
Som i vissa sekter är det möjligt att döda en process om du vet dess rätta namn.
		-- Ken Thompson and Dennis M. Ritchie

%
Som i protestantiska Europa, däremot, där sekter delas oändligt inmindre konkurrerande sekter och ingen kyrka dominerade alla andra, är alla olikai den fragmenterade värld IBM. Det området är nu ett kaos av motstridiganormer och standarder som inte ens IBM kan hoppas på att styra. Du kan köpa endator som fungerar som en IBM-maskin, men innehåller ingenting görs eller säljs avIBM själv. Renegades från IBM ständigt ställa upp konkurrerande företag och inrättastandarderna för deras egen. När IBM övergav nyligen en del av sin ursprungligastandarder och förordnas nya, många av sina konkurrenter förklarade en puritantrohet till IBM: s ursprungliga tro, och fördömde företaget som en splittrandeinnovatör. Ändå är IBM världen förenas av sin misstro mot ikoner ochbilder. IBM: s skärmar är utformade för språket, inte bilder. GravenBilderna kan tolereras av de lyxiga kulter, men den sanna IBM tron ​​förlitarpå åtstramning av ordet.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Så länge som det finns dåligt definierade mål, bisarra buggar och orealistiskscheman, kommer det att finnas Real Programmerare villiga att hoppa in och lösaProblemet, spara dokumentation för senare.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Från och med nästa torsdag, kommer UNIX spolas till förmån för TOPS-10.Uppdatera dina program.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Från och med nästa tisdag, kommer C spolas till förmån för COBOL.Uppdatera dina program.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Från och med nästa vecka kommer lösenord föras in i morsekod.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Som en del av ett pågående arbete för att hålla dig, Fortune läsare, à jour medden värdefull information som dagligen korsar Usenet, Fortune presenterar:Nyhetsartiklar som svarar * dina * frågor, # 1:Nyhetsgrupper: comp.sources.dÄmne: Hur gör jag kör C-kod som tas emot från källorNyckelord: C källorDistribution: naJag vet inte hur man ska köra C-program som läggs ikällor diskussionsgrupp. Jag spara filerna, redigera dem för att ta bortrubriker och ändra läge så att de är körbara, men jagkan inte få dem att köra. (Jag har aldrig skrivit ett C-program tidigare.)De måste sammanställas? Med vilken kompilator? Hur gör jag? OmJag sammanställa dem, är ett objektkoden fil som genereras eller måste jag skapauttryckligen med> karaktär? Finns det något annat som	måste göras?
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Som en del av omvandlingen, dataspecialister skrev 1500 program;en process som traditionellt kräver viss felsökning.omvandling till ett nytt datasystem.
		-- USA Today, referring to the Internal Revenue Service

%
Så snart vi började programmering, fann vi till vår förvåning att det inte varså lätt att få program direkt som vi hade trott. Debugging var tvungen att varaupptäckt. Jag kommer ihåg den exakta ögonblick när jag insåg att en stordel av mitt liv därefter skulle spenderas i att hitta fel imina egna program.
		-- Maurice Wilkes, designer of EDSAC, on programming, 1949

%
Eftersom systemet kommer upp, kommer komponentbyggare från tid till annan visasbärande heta nya versioner av sina pjäser - snabbare, mindre, mer kompletta,eller förmodat mindre buggy. Ersättandet av en arbetande komponent med en nyversionen kräver samma systematiska testförfarande som lägger till en nykomponent gör, även om det skulle kräva mindre tid för mer komplett ocheffektiva testfall vanligtvis tillgängliga.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Som livets prövningar fortsätter att ta sin tribut, kom ihåg att detär alltid en framtid i adb.
		-- National Lampoon, "Deteriorata"

%
Som Will Rogers skulle ha sagt, "Det finns inget sådant som en gratis variabel."
		-- National Lampoon, "Deteriorata"

%
ASCII en dum fråga, får du en EBCDIC svar.
		-- National Lampoon, "Deteriorata"

%
Aska, DOS till DOS.
		-- National Lampoon, "Deteriorata"

%
Fråga inte för vem <CONTROL-G> vägtullar.
		-- National Lampoon, "Deteriorata"

%
Assembler erfarenhet är [viktigt] för löptidenoch förståelse för hur datorer fungerar som det ger.
		-- D. Gries

%
Asynkrona ingångar är roten till våra ras problem.
		-- D. Winker and F. Prosser

%
Vid ungefär 2500 e Kr, upptäcker mänskligheten ett datorproblem som * måste * varalöst. Den enda svårigheten är att problemet är NP-fullständig och viljata tusentals år även med den senaste optiska biologiska tekniktillgängliga. De bästa datavetare sitta ner för att tänka ut någon lösning.I stor bestörtning, en av C.S. folk berättar man om det. Detär bara en lösning, säger han. Kom ihåg fysik 103, modern fysik, allmänrelativitet och alla. Hon svarar: "Vad har det att göra med att lösaett datorproblem? ""Kom ihåg det dubbla paradox?"Efter några minuter, säger hon, "jag skulle kunna sätta datorn på en mycketsnabb maskin och datorn skulle ha bara ett par minuter att beräkna mensom är raka motsatsen till vad vi vill ... Självklart! Lämnadator här, och påskynda jorden! "Problemet var så viktigt att de gjorde precis det. Närjorden kom tillbaka, de presenteras med svaret:IEH032 Fel i JOBB styrkortet.
		-- D. Winker and F. Prosser

%
Vid en första anblick är idén om några regler eller principer överlagras pådet kreativa sinnet verkar mer troligt att hindra än att hjälpa, men det ärganska osann i praktiken. Disciplinerat tänkande fokuserar inspiration snarareän blinkers den.
		-- G. L. Glegg, "The Design of Design"

%
På koncernnivå L, Stoffel övervakar sex första klassens programmerare, en ledandeutmana ungefär jämförbar med vallning katter.
		-- The Washington Post Magazine, 9 June, 1985

%
Vid källan varje fel som skylls på datorn hittar duåtminstone två mänskliga fel, inklusive felet att skylla det på datorn.
		-- The Washington Post Magazine, 9 June, 1985

%
Undvik konstiga kvinnor och tillfälliga variabler.
		-- The Washington Post Magazine, 9 June, 1985

%
Basic är en hög nivå languish. APL är en hög nivå ångest.
		-- The Washington Post Magazine, 9 June, 1985

%
BASIC är datavetenskap motsvarande `vetenskaplig kreationism".
		-- The Washington Post Magazine, 9 June, 1985

%
BASIC är att datorprogrammering som QWERTY är att skriva.
		-- Seymour Papert

%
Var försiktig när en slinga lämnar till samma plats från sidan och botten.
		-- Seymour Papert

%
Bakom varje stor dator sitter en mager liten nörd.
		-- Seymour Papert

%
Bell Labs Unix - Nå ut och grep någon.
		-- Seymour Papert

%
Akta dig för buggar i ovanstående kod; Jag har bara visat det riktigt, inte provat det.
		-- Donald Knuth

%
Akta dig för Programmerare som bär skruvmejslar.
		-- Leonard Brandwein

%
Akta dig för Turing Tar-grop där allt är möjligt, men inget avintresse är lätt.
		-- Leonard Brandwein

%
Akta nya TTY-koden!
		-- Leonard Brandwein

%
Blinding hastighet kan kompensera för en hel del brister.
		-- David Nichols

%
Båda modellerna är identiska i prestanda, funktionell drift, ochgränssnitt kretsdetaljer. De två modellerna, dock är inte kompatiblapå samma kommunikationsledning anslutning.
		-- Bell System Technical Reference

%
Håll i er. Vi är på väg att prova något som gränsar till det unika:en faktiskt ganska allvarlig teknisk bok som inte bara (gasp) häftigtanti-Solemn, men också (rysning) tar sidor. Jag brukar tänka på det som`Konstruktiv Snottiness."
		-- Mike Padlipsky, "Elements of Networking Style"

%
Hjärna stekt - Kärna dumpas
		-- Mike Padlipsky, "Elements of Networking Style"

%
Bredd-först-sökning är bulldozer vetenskap.
		-- Randy Goebel

%
Brian Kernighan har en bil som han hjälpte design.Till skillnad från de flesta bilar har varken hastighetsmätare eller gas mätare, ellernågon av de många idiot lampor som plågar den moderna föraren.Snarare om föraren gör några misstag, en jätte "?" lyser imitten av instrumentbrädan. "Den erfarna förare", säger han, "kommeroftast vet vad som är fel. "
		-- Randy Goebel

%
Föra datorer i hemmet kommer inte att ändra något av det, men kanvitalisera hörnet salong.
		-- Randy Goebel

%
Bygga ett system som även en dåre kan använda och bara en idiot kommer att vilja använda den.
		-- Randy Goebel

%
Att bygga översättare är bra rent nöje.
		-- T. Cheatham

%
Bussfel - drivrutin utförs.
		-- T. Cheatham

%
Bussfel - lämna den bakre luckan.
		-- T. Cheatham

%
Men i vår entusiasm, kunde vi inte motstå en radikal översyn avsystem där alla dess stora brister har varit utsatt,analyseras, och ersätts med nya svagheter.
		-- Bruce Leverett, "Register Allocation in Optimizing Compilers"

%
Men det har tagit oss långt bort från gränssnittet, vilket inte är en dåligplats att vara, eftersom jag särskilt vill gå vidare till kludge.Varför människor har så mycket problem att förstå kludge? Vadär en kludge, trots allt, men inte tillräckligt K: s, inte tillräckligt ROM, intetillräckligt RAM, dålig kvalitet gränssnitt och för få byte för att gå runt?Har jag förklarade ännu om byte?
		-- Bruce Leverett, "Register Allocation in Optimizing Compilers"

%
"Men vad vi behöver veta är, gör människor vill nasalt inför datorer?"
		-- Bruce Leverett, "Register Allocation in Optimizing Compilers"

%
Genom lång tradition, jag tar tillfället i akt stund andradesigners i tunn förklädnad av god, ren kul.Fool kolumn.
		-- P. J. Plauger, "Computer Language", 1988, April

%
BYTE redaktörer är människor som skiljer agnarna från vetet, och sedanförsiktigt ut vetet.
		-- P. J. Plauger, "Computer Language", 1988, April

%
Byte tungan.
		-- P. J. Plauger, "Computer Language", 1988, April

%
C-koden.C Code Kör.Kör, kod, KÖR!	SNÄLLA DU!!!!
		-- P. J. Plauger, "Computer Language", 1988, April

%
C själv.
		-- P. J. Plauger, "Computer Language", 1988, April

%
C gör det enkelt för dig att skjuta dig själv i foten. C ++ gör atthårdare, men när du gör, blåser det bort hela benet.
		-- Bjarne Stroustrup

%
C'est magnifique, mais ce n'est pas l'Informatique.
		-- Bosquet [on seeing the IBM 4341]

%
C ++ är det bästa exemplet på andra systemet effekt, eftersom OS / 360.
		-- Bosquet [on seeing the IBM 4341]

%
... C ++ erbjuder ännu mer flexibel kontroll över synlighet medlemobjekt och medlemsfunktioner. Specifikt kan medlemmar placeras ioffentliga, privata eller skyddade delar av en klass. Medlemmar deklareras ioffentliga delar är synliga för alla kunder; medlemmar förklarade i den privatadelar är helt inkapslade; och medlemmar deklareras i de skyddade delarnaär synliga endast till själva klassen och dess underklasser. C ++ stöder ocksåbegreppet * _______ vänner *: kooperativa klasser som har tillåtelse att se varjeandra privata delar.
		-- Grady Booch, "Object Oriented Design with Applications"

%
Lugna ner, är det * ____ bara * ettor och nollor.
		-- Grady Booch, "Object Oriented Design with Applications"

%
Det går inte att öppna / usr / share / games / förmögenheter / förmögenheter. Lock fastnat på kakburken.
		-- Grady Booch, "Object Oriented Design with Applications"

%
Kan inte öppna /usr/share/games/fortunes/fortunes.dat.
		-- Grady Booch, "Object Oriented Design with Applications"

%
CChheecckk yyoouurr dduupplleexx sswwiittcchh ..
		-- Grady Booch, "Object Oriented Design with Applications"

%
CCI Ström 6/40: en styrelse, en megabyte cache och en attityd ...
		-- Grady Booch, "Object Oriented Design with Applications"

%
Center möte på 4:00 i 2C-543.
		-- Grady Booch, "Object Oriented Design with Applications"

%
Civilisation, som vi känner den, kommer att sluta någon gång denna kväll.Se SYSNOTE morgon för mer information.
		-- Grady Booch, "Object Oriented Design with Applications"

%
COBOL är för morons.
		-- E. W. Dijkstra

%
Cobol programmerare är deppig.
		-- E. W. Dijkstra

%
Kodning är lätt; Allt du behöver göra är att sitta stirrar på en terminal tills dropparnablod formulär på din panna.
		-- E. W. Dijkstra

%
Jämföra software engineering klassisk teknik förutsätter att programvarahar förmågan att bära ut. Programvaran fungerar normalt, eller inte. Detantingen fungerar eller inte. Programvara i allmänhet inte försämra, slipa,stretch, twist, eller avlägsna. Att behandla det som en fysisk enhet, därför ärfelaktig tillämpning av våra ingenjörskunskaper. Klassiska ingenjörs behandlaregenskaperna av hårdvara; programvaruteknik bör ta itu medegenskaper * programvara *, och inte med hårdvara eller ledning.
		-- Dan Klein

%
KOMPASS [för CDC-6000-serien] är den typ av assembler man förväntar sig avett företag vars president koder oktala.
		-- J. N. Gray

%
... Hårdvara framsteg är så snabb. Ingen annan teknik sedancivilisation började har sett sex storleksordningar i prestations prisvinna på 30 år.
		-- Fred Brooks

%
Programmerare gör det byte av byte.
		-- Fred Brooks

%
Programmerare dör aldrig, de bara gå vilse i behandlingen.
		-- Fred Brooks

%
Datorprogram expandera för att fylla kärnan tillgänglig.
		-- Fred Brooks

%
Datavetenskap är enbart efter Turing nedgång i formella systemteori.
		-- Fred Brooks

%
Computer Science är den enda disciplin där vi ser att lägga till en ny flygeltill en byggnad som underhåll
		-- Jim Horning

%
Datorer är inte intelligent. De tror bara de är.
		-- Jim Horning

%
Datorer är opålitliga, men människor är ännu mer opålitliga.Varje system som beror på mänsklig tillförlitlighet är opålitlig.
		-- Gilb

%
Datorer är värdelösa. De kan bara ge dig svar.
		-- Pablo Picasso

%
Datorer kan räkna ut alla typer av problem, förutom de saker ivärlden som bara inte lägga upp.
		-- Pablo Picasso

%
Datorer egentligen inte tänka.Du tror bara att de tror.		(Vi tror.)
		-- Pablo Picasso

%
Datorer kommer inte att fulländade tills de kan räkna ut hur mycket merän uppskattningen jobbet kommer att kosta.
		-- Pablo Picasso

%
Begrepps integritet i sin tur kräver att konstruktionen måste fortsättafrån ett sinne, eller från ett mycket litet antal enas resonans sinnen.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
grattis! Du är den miljonte användare att logga in i vårt system.Om det finns något speciellt vi kan göra för dig, vad som helst, intetveka att fråga!
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Cosmotronic Software Obegränsad Inc. garanterar inte attfunktionerna i programmet uppfyller dina krav eller attdriften av programmet kommer att vara oavbruten eller felfri.Men Cosmotronic Software Unlimited Inc. motiverardiskett (er) på vilken programmet är inredda för att vara svart färg ochkvadratisk form vid normal användning under en period av nittio (90) dagar fråninköpsdatum.OBS: UNDER INGA OMSTÄNDIGHETER COSMOTRONIC SOFTWARE UNLIMITED ELLERDistributörer och deras ÅTERFÖRSÄLJARE VARA ANSVARIGA FÖR NÅGRA SKADOR, INKLUSIVENÅGON FÖRLUST AV VINST, FÖRLORADE BESPARINGAR, förlorade tålamodet ELLER ANNAN TILLFÄLLIG ELLERSKADOR.
		-- Horstmann Software Design, the "ChiWriter" user manual

%
Det gick inte att vi jury-rig katten att fungera som en ljud switch, och har det skrikapå människor att spara sina kärn bilder innan du loggar ut dem? jag är säkerprod boskap skulle vara effektivt i detta avseende. I varje fall, en traversmonterad leguan, medan mer perversa, ger bättre dragkraft, för att inte tala omär lättare att satsa.
		-- Horstmann Software Design, the "ChiWriter" user manual

%
Räkna i binärt är precis som att räkna i decimal - om du är alla tummar.
		-- Glaser and Way

%
Räkna i oktala är precis som att räkna i decimal - om du inte använder tummarna.
		-- Tom Lehrer

%
[Crash program] misslyckas eftersom de är baserade på teorin att, med niokvinnor gravida, kan du få en baby i månaden.
		-- Wernher von Braun

%
Crazee Edeee hans priserna är galen !!!
		-- Wernher von Braun

%
Att skapa datorprogram är alltid en krävande och mödosamtprocess - en övning i logik, tydligt uttryck, och nästan fanatiskuppmärksamhet på detaljer. Det kräver intelligens, engagemang och enenormt hårt arbete. Men en viss oförutsägbaroch ofta unrepeatable inspiration är det som gör vanligtvis skillnadenmellan tillräcklighet och kvalitet.
		-- Wernher von Braun

%
VMS-F-PDGERS, pudding mellan öronen
		-- Wernher von Braun

%
Kära Emily, hur testmeddelanden?Kära berörs:Det är viktigt, när man testar, för att testa hela nätet. aldrig testetbara ett subnät fördelning när hela nätet kan göras. Också sätta "vänligenignorera "på dina testmeddelanden, eftersom vi alla vet att alla alltid hopparett meddelande med en rad liknande. Använd inte ett ämne som "mitt kön är kvinnligtmen jag kräver att behandlas som män. "eftersom sådana artiklar läses på djupetav alla USEnauts.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Hur kan jag välja vilka grupper för att skriva in?Kära förvirrad:Plocka så många som möjligt, så att du får en bred publik. Efterallt finns på nätet för att ge dig en publik. Ignorera dem som föreslår att dubör endast använda grupper där du tror att artikeln är mycket lämpligt.Välj alla grupper där vem som helst kan även vara lite intresserad.Se alltid till uppföljningar gå till alla grupper. I de sällsynta fallatt du lägger en uppföljning som innehåller något originellt, se till att duutöka listan över grupper. Aldrig innehålla en "Uppföljning till:" linje iheader, eftersom vissa människor kan missa en del av den värdefulla diskussionde marginella grupper.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Jag samlade svar på en artikel jag skrev, och nu är det dags attsammanfatta. Vad ska jag göra?Kära redaktör:Helt enkelt slå samman alla artiklar ihop till en stor fil och postden där. På Usenet, kallas detta en sammanfattning. Det låter folk läsa allasvar utan irriterande nyhetsläsare i vägen. Gör samma sak närsammanfattar en röst.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Jag läste nyligen en artikel som sa, "svara per post, jag ska sammanfatta."Vad ska jag göra?Dear Tveksamt:Lägg upp ditt svar till hela nätet. Denna begäran gäller endastdumma människor som inte har något intressant att säga. Dina inlägg ärmycket mer lönsamt än andra folk, så det skulle vara ett slöseri att svara genombrev.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Jag såg en lång artikel som jag vill motbevisa noga, vad skaJag gör?Kära Arg:Inkludera hela texten med din artikel, och inkludera dina kommentarermellan raderna. Var noga med att göra det och inte skicka, även om din artikelser ut som ett svar till den ursprungliga. Alla * älskar * att läsa de långapunkt för punkt debatter, särskilt när de utvecklas till utskällningar ochmassor av "Är också!" -- "Är inte!" - "Är för, twizot!" utbyten.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Jag har allvarliga meningsskiljaktigheter med någon på nätet. jagförsökte klagomål till hans sysadmin, organisera postkampanjer, som kallas förhans avlägsnande från nätet och ringa sin arbetsgivare för att få honom sparken.Alla skrattade åt mig. Vad kan jag göra?Kära berörs:Gå till dagstidningar. De flesta moderna reportrar är top-notch datorexperter som förstår nätet, och dina problem, perfekt. Deskriver ut noggranna, motiverade berättelser utan några fel alls, och säkertrepresenterar situationen korrekt för allmänheten. Allmänheten kommer också allahandla klokt, eftersom de är också fullt medveten om de subtila natur nettosamhälle.Papper aldrig sensation eller snedvrida, så se till att påpeka sakersom rasism och sexism varhelst de kan finnas. Var noga samt att deförstå att allt på nätet, särskilt förolämpningar, menasbokstavligen. Länk vad som framkommer på nätet för att orsakerna till Förintelsen, ommöjlig. Om vanliga papper inte kommer att ta historien, gå till en tabloid papper -de är alltid intresserade av bra historier.Genom att arrangera allt detta gratis publicitet för nätet, kommer du att bli mycketvälkända. Människor på nätet kommer att vänta i spänd förväntan för varjebokföring, och hänvisar till dig hela tiden. Du får mer post än du någonsintrodde var möjligt - den ultimata netto framgång.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Jag är fortfarande förvirrad om vilka grupper artiklar ska bokförastill. Vad sägs om ett exempel?Käre Still:Ok. Låt oss säga att du vill rapportera att Gretzky har handlats frånOilers till Kings. Nu genast du kanske tror rec.sport.hockeyskulle vara tillräckligt. FEL. Många fler människor kan vara intresserade. Det här är enstor handel! Eftersom det är en nyhetsartikel, hör det i nyheterna. * Hierarkinockså. Om du är en nyhets admin, eller om det finns en på din dator, försöknews.admin. Om inte, använd news.misc.De Oilers är förmodligen intresserad av geologi, så försök sci.physics.Han är en stor stjärna, så post till sci.astro och sci.space eftersom de är ocksåintresserad av stjärnor. Därefter är hans namn polska klingande. Så skicka tillsoc.culture.polish. Men den gruppen inte existerar, så kors post tillnews.groups tyder det bör skapas. Med så här många grupper avintresse, kommer din artikel vara ganska bisarra, så skicka till talk.bizarre somväl. (Och lägga till comp.std.mumps, eftersom de knappast få några artiklardär, och en "comp" grupp kommer att fortplanta din artikel ytterligare.)Du kan också finna det är roligare att skriva artikeln en gång i varjegrupp. Om du lista alla diskussionsgrupper i samma artikel, några diskussionsgruppsläsareendast visa artikeln till läsaren en gång! Inte tolerera detta.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Emily:Idag har jag skrivit en artikel och glömde att inkludera min signatur.Vad ska jag göra?Dear Glömsk:Rusa till din terminal direkt och skickar en artikel som säger,"Oj, jag glömde att lägga min signatur med den sista artikeln. Härdet är."Eftersom de flesta människor kommer att ha glömt tidigare artikel,(Särskilt eftersom det vågade vara så tråkigt att inte ha en trevlig, saftigsignatur) Detta kommer att påminna dem om det. Dessutom människor bryr sig mycket merom signaturen i alla fall.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Käre Ms Postnews:Jag kunde inte få e-post fram till någon på en annan plats. Vad	borde jag?Kära Eager:Inga problem, bara skicka ditt meddelande till en grupp som många människorläsa. Säg, "Detta är för John Smith. Jag kunde inte få e-post via så jag ärlägga ut den. Alla andra vänligen ignorera. "På detta sätt tiotusentals människor kommer att spendera några sekunder scanningöver och ignorerar din artikel, med upp över 16 mantimmar deras kollektivatid, men du kommer att sparas den fruktansvärda problem att kontrollera genom usenetkartor eller letar efter alternativa rutter. Tänk om du inte kunde fördeladitt meddelande till 9000 andra datorer, kan du faktiskt behöva (gasp) samtalnummerupplysningen för 60 cent, eller ens ringa person. Detta kan kostaså mycket som några dollar (!) för en 5 minuters samtal!Och visst är det bättre att spendera 10 till 20 dollar i andraspengar att fördela meddelandet än för dig att ha att slösa $ 9 på en övernattningbrev, eller till och med 25 cent på ett frimärke!Glöm inte. Världen kommer att upphöra om ditt meddelande inte komma igenom,så skicka det så många platser som möjligt.
		-- Emily Postnews Answers Your Questions on Netiquette

%
Dear Sir,Jag motsätter sig spridning av mikrochips antingen till hemmet ellertill kontoret, har vi mer än nog av dem prackas på oss offentligtplatser. De är en motbjudande amerikanism, och kan bara resultera i böndernatvingas att växa mindre potatis, vilket i sin tur kommer att leda till massiv oföranställning i den redan allvarligt deprimerad jordbruksindustrin.Med vänlig hälsning,Capt. Quinton D'Arcy, J.P.Seven
		-- Letters To The Editor, The Times of London

%
Debug är mänsklig, de-fix gudomlig.
		-- Letters To The Editor, The Times of London

%
DEC diagnostik skulle köras på en död val.
		-- Mel Ferentz

%
#define BITCOUNT (x) (((BX_ (x) + (BX_ (x) >> 4)) & 0x0F0F0F0F)% 255)#define BX_ (x) ((x) - (((x) >> 1) & 0x77777777) \- (((X) >> 2) & 0x33333333) \- (((X) >> 3) & 0x11111111))
		-- really weird C code to count the number of bits in a word

%
(Defun NF (a c)  (Dir ((null c) ())((Atom (bil c))(Bifoga (lista (eval (lista 'getchar (lista (bil c) a) (CADR c))))(Nf en (cddr c))))(T (bifoga (lista (imploderar (nf en (bil c)))) (nf en (CDR c))))))(Defun AD (vill arbetsplatsen utmana Boston-området)  (cond   ((Eller (ej (lika vill-jobb "ja))(Inte (lika boston-område "ja))(Lessp utmanande 7)) ())   (T (bifoga (nf (få "ad" expr)((Caaddr en caadr två bil en bil 1)(Bil 5 cadadr 9 cadadr 8 cadadr 9 caadr 4 bil 2 bil 1)(Bil 2 caadr 4)))      (Lista "851-5071x2661)))));;; Vi är en positiv särbehandling arbetsgivare.
		-- really weird C code to count the number of bits in a word

%
Leverera igår, kod idag, tror morgon.
		-- really weird C code to count the number of bits in a word

%
Visste du att för priset av en 280-Z kan du köpa två Z-80-talet?
		-- P. J. Plauger

%
Olika all krånglig en av i labyrinten är du, passager lite.
		-- P. J. Plauger

%
Digitala kretsar tillverkas från analoga delar.
		-- Don Vonada

%
Diskutrymme - finalgränsen!
		-- Don Vonada

%
DISCLAIMER:Användning av denna avancerade datortekniken innebär inte ett godkännandeVäst industriella civilisationen.
		-- Don Vonada

%
Varning: "Dessa yttranden är mina egna, men för en liten avgift de varadin också."
		-- Dave Haynie

%
Disk kris, vänligen städa upp!
		-- Dave Haynie

%
Diskar resa i förpackningar.
		-- Dave Haynie

%
Disraeli var ganska nära: faktiskt finns Lies, Damn lögner, statistik,Riktmärken och leveransdatum.
		-- Dave Haynie

%
Inte lägga sig i angelägenheter troff, för det är subtil och snar till vrede.
		-- Dave Haynie

%
Inte förenkla utformningen av ett program om kan hittat ett sätt att göradet komplexa och underbart.
		-- Dave Haynie

%
Använd inte de blå knapparna på denna terminal.
		-- Dave Haynie

%
Vet ni vad du gör, eller är du bara hacka?
		-- Dave Haynie

%
*** HAR NI en rastlös lust att programmet? ***Vill du omedelbar respekt som kommer från att kunna använda teknisktermer som ingen förstår? Vill du sätta skräck och avsky ihjärtan DP chefer överallt? Om så är fallet, låt den berömda programmerare "Skola leda dig på ... i en värld av professionell datorprogrammering.*** Programmerar FÖR DIG? ***Programmering är inte för alla. Men om du har lust att lära, vi kanhjälpa dig att komma igång. Allt du behöver är den berömda programmerare "Course ochtillräckligt med pengar för att hålla dessa lektioner kommer månad efter månad.*** Ta vår gratis Högskoleprov ***För att avgöra om du är kvalificerad att vara en programmerare, ta en stund attprova detta enkla test:(1) Skriv ner siffrorna noll till nio och de första sex bokstäveri alfabetet (Tips: 0123456789ABCDEF).(2) vars bild finns på baksidan av en tjugodollarsedel?(3) Vad är statens huvudstad Idaho?Om du lyckats läsa alla tre frågor utan att undra varför vi frågadedem, kan du ha en framtid som programmerare.
		-- Dave Haynie

%
Lider du smärtsam eliminering?Lider du smärtsam recrimination?Lider du smärtsam belysning?Lider du smärtsam hallucination?
		-- Don Juan, cited by Carlos Casteneda

%
Dokumentation är som sex: när det är bra, det är mycket, mycket bra; ochnär det är dåligt, är det bättre än ingenting.
		-- Dick Brandon

%
Dokumentation är ricinolja programmering.Chefer vet att det måste vara bra eftersom de programmerare hatar det så mycket.
		-- Dick Brandon

%
Har en bra bonde försummar en gröda han har planterat?Har en bra lärare förbise även de mest ödmjuka student?Har en god far låta ett enda barn att svälta?Har en bra programmerare vägra att behålla sin kod?
		-- Geoffrey James, "The Tao of Programming"

%
Jämför inte flyttal enbart för jämställdhet.
		-- Geoffrey James, "The Tao of Programming"

%
Bli inte lurade in av kommentarerna - de kan vara fruktansvärt missvisande.Debug bara kod.
		-- Dave Storer

%
Inte slår an tangenterna så hårt, det gör ont.
		-- Dave Storer

%
Inte svettas det - det är bara ettor och nollor.
		-- P. Skelly

%
DOS Air:Alla passagerare går ut på landningsbanan, greppa tag i planet, driva dettills det blir i luften, hoppa på, hoppa av när den träffar marken igen.Sedan ta tag i planet igen, skjut tillbaka den i luften, hoppa på etcetera.
		-- P. Skelly

%
DOS öl: kräver att du använder din egen konservöppnare, och kräver att duLäs instruktionerna noga innan du öppnar burken. ursprungligen barakom i en 8-oz. kan, men nu kommer i en 16-oz. Kan. Emellertid är burkindelat i 8 fack i 2 oz. vardera, vilket måste nåsseparat. Snart ska avbrytas, även om en hel del människor kommeratt hålla dricka det efter att det inte längre är tillgänglig.
		-- P. Skelly

%
På grund av brist på diskutrymme, har denna förmögenhet databas avbrutits.
		-- P. Skelly

%
Under de följande två timmarna, kommer systemet att gå upp och ned fleragånger, ofta med lin ~ Po '~ {po ~ poz ~ PPO \ ~ {på ~ Po' ~ {o [po ~ y oodsou> # w4k ** n ~ Po '~ {ol; lkld, f, g, dd; po \ ~ {o
		-- P. Skelly

%
E Pluribus Unix
		-- P. Skelly

%
Varje ny användare av ett nytt system avslöjar en ny klass av buggar.
		-- Kernighan

%
Var och en av dessa sekter motsvarar en av de två antagonisterna i en ålder avReformation. I sfären av Apple Macintosh, som i katolska Europa,tillbedjare inbördes andäktigt in skärmar fyllda med "ikoner". Allt är sund ochbilder och Appledom. Även ord ser ut som dekorativa filigrees i exotiskatypsnitt. Den största ikonen för alla, okränkbara Apple själva, står iden dominerande position vid det övre vänstra hörnet av skärmen. En centralhuvudkontor påbjuder form av alla riter och praxis.Infalliable läran frågor från en verkställande tjänsteman vars urval skeri ett förseglat styrelserum. Skulle någon i hans curia ifrågasätta hans befogenheter,gärningsmannen är bannlyst i mörkret. Det utdrivna kättare grundarett nytt bolag, muttrar dunkelt av den kommande ålder och nästa gång datorn,sedan försvinner in i tystnad, med hans eget med honom. MammanFöretaget förbjuder finansiella konkurrens strängt som den kväver ideologiskkonkurrens; Om du vill använda datorprogram som följer Applesortodoxi, måste du köpa en dator tillverkas och säljs av Apple själva.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
/ Jorden är 98% full ... du ta bort någon du kan.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Jorden är en beta webbplats.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
/ Jorden filsystem fullt.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Einstein menade att det måste förenklas förklaringar av naturen, eftersomGud är inte nyckfull eller godtycklig. Ingen sådan tro tröstar programvaraningenjör.
		-- Fred Brooks

%
Lika byte för kvinnor.
		-- Fred Brooks

%
Fel i operatör: lägg öl
		-- Fred Brooks

%
Etablerad teknik tenderar att kvarstå i ansiktet av ny teknik.
		-- G. Blaauw, one of the designers of System 360

%
Eudaemonic forskning fortsatte med den avslappnade mani utmärkande för denna del avvärlden. Naken sola på baksidan däck kombinerades med telefonsamtal tillAvancerade Kinetics i Costa Mesa, American Laser Systems i Goleta, AutomationIndustries i Danbury, Connecticut, Arenberg Ultraljud i Jamaica Plain,Massachusetts, och Hewlett Packard i Sunnyvale, Kalifornien, där NormanPackards kusin, David, som ordförande i styrelsen. Tricket var attgöra dessa samtal vid middagstid, i hopp om att ut-till-lunch chefer skulle återvändadem på egen bekostnad. Eudaemonic Enterprises, för alla de visste, kanskeen snabbväxande dataföretag förgrening av Silicon Valley. sniffningmöjligheten till hög volym försäljning, dessa chefer lite misstänkt attde talade på den andra änden av linjen till en naken fysiker galenöver roulette.
		-- Thomas Bass, "The Eudaemonic Pie"

%
<<<<< Utrymningsväg <<<<<
		-- Thomas Bass, "The Eudaemonic Pie"

%
Även byte får ensam för lite.
		-- Thomas Bass, "The Eudaemonic Pie"

%
Någonsin undrat om ursprunget till begreppet "buggar" som tillämpas på datornteknologi? US Navy Capt. Grace Murray Hopper har förstahands förklaring.74-årige kaptenen, som fortfarande är i aktiv tjänst, var en pionjär inomdatateknik under andra världskriget. Vid CW Post Center of LongIsland University, Hopper berättade en grupp av Long Island kommunal skola administrativamännen att den första datorn "bug" var en riktig bugg - en mal. vid Harvarden augustinatt 1945, var Hopper och hennes medarbetare som arbetar på"Morfar" av moderna datorer, var Mark I. "Saker går dåligt;det var något fel i en av kretsarna i den långa inglasadedator ", sade hon." Slutligen, någon hittat oroshärd och med hjälp avvanliga pincett, bort problemet, en två-tums mal. Från och med då, närnågot gick fel med en dator, sa vi att det hade fel i det. "Hoppersade att när sanningshalten i hennes berättelse ifrågasattes nyligen, "jag hänvisadedem till min 1945 loggbok, nu i samlingen av Naval Surface VapenCenter, och de fann resterna av det mal tejpade till sidan ifråga."[Faktiskt termen "bug" hade ännu tidigare användning ibeaktande av problem med radio hårdvara. Ed.]
		-- Thomas Bass, "The Eudaemonic Pie"

%
"Varje grupp har ett par experter. Och varje grupp har åtminstone enidiot. Således är balans och harmoni (och oenighet) upprätthålls. Dessibland svårt att komma ihåg detta i huvuddelen av de e-gräl som allaav krångel och smärta orsakas vanligtvis av en eller två högt motiverade,kaustiska twits. "
		-- Chuq Von Rospach, about Usenet

%
Varje program har åtminstone en bug och kan förkortas genom åtminstone ettinstruktion - från vilken genom induktion, kan man dra slutsatsen att varjeProgrammet kan reduceras till en instruktion som inte fungerar.
		-- Chuq Von Rospach, about Usenet

%
Varje program är en del av något annat program, och sällan passar.
		-- Chuq Von Rospach, about Usenet

%
Varje Solidaritet center hade högar och högar av papper ... alla varäter papper och en polis var vid dörren. Allt du behöver göra är attböja en disk.kommenterade fördelarna med att använda datorer i stödav deras rörelse.
		-- A member of the outlawed Polish trade union, Solidarity,

%
Alla behöver lite kärlek någon gång; sluta hacka och förälska!
		-- A member of the outlawed Polish trade union, Solidarity,

%
Alla kan lära sig att skulptera: Michelangelo skulle ha behövt varalära ___ inte. Så är det med de stora programmerare.
		-- A member of the outlawed Polish trade union, Solidarity,

%
Evolution är en miljon linje datorprogram faller på plats av en slump.
		-- A member of the outlawed Polish trade union, Solidarity,

%
Överdriven inloggning eller utloggning meddelanden är ett säkert tecken på senilitet.
		-- A member of the outlawed Polish trade union, Solidarity,

%
ANLÄGGNING godtas 100044200000;
		-- A member of the outlawed Polish trade union, Solidarity,

%
Känsla amorös, såg hon under bladen och ropade: "Åh, nej,Det är Microsoft! "
		-- A member of the outlawed Polish trade union, Solidarity,

%
Fellow programmerare, hälsningar! Du läser ett brev som kommer att föradu tur och lycka. Bara post (eller UUCP) tio kopior av detta brevtill tio av dina vänner. Innan du gör kopior, skicka ett chip ellerannan bit av hårdvara, och 100 rader C-kod till den första personen pålista ges längst ner i detta brev. Sedan ta bort deras namn och lägga tiller till botten av listan.Bryt inte kedjan! Gör kopian inom 48 timmar. Gerald R. från SanDiego misslyckats med att sända ut sina tio exemplar och vaknade nästa morgon att hittahans arbetsbeskrivning ändras till "COBOL programmerare." Fred A. New York skickasut sina tio exemplar och inom en månad hade nog hårdvara och mjukvara för attbygga en Cray tillägnad spela Zork. Martha H. från Chicago skrattade åtdetta brev och bröt kedjan. Kort därefter utbröt en brand ihennes terminal och hon tillbringar nu sina dagar skriva dokumentation för IBM PC.Bryt inte kedjan! Skicka ut dina tio exemplar idag!
		-- A member of the outlawed Polish trade union, Solidarity,

%
Till exempel, om \ thinmskip = 3mu, detta gör \ thickmskip = 6mu. Men omdu också vill använda \ skip12 för horisontell lim, vare sig i matematikläge ellerinte, kommer mängden hoppa vara i punkter (t ex 6pt). Regeln äratt lim i matematikläge varierar med storleken endast när det är en \ mskip;när du flyttar mellan ett mskip och vanlig hoppa över, omräkningsfaktorn1mu = 1pt används alltid. Innebörden av "\ mskip \ skip12" och'\ Baselineskip = \ den \ thickmskip "ska vara klar.
		-- Donald Knuth, TeX 82 -- Comparison with TeX80

%
Fly Windows NT:Alla passagerare utför sina platser ut på asfalten, placera stolarnai konturerna av en plan. Alla sitter ner, flaxa med armarna och göra jetswooshing låter som om de flyger.
		-- Donald Knuth, TeX 82 -- Comparison with TeX80

%
"För övrigt, jämföra din fickdator med de massiva jobbtusen år sedan. Varför inte då det sista steget för att göra sig av meddatorer helt och hållet? "
		-- Jehan Shuman

%
FORTH IF TUTA DÅ
		-- Jehan Shuman

%
FORTRAN är ett bra exempel på ett språk som är lättare att tolkamed hjälp av ad hoc-tekniker.[Vad är bra om det? Ed.]
		-- D. Gries

%
FORTRAN är inte en blomma, men ett ogräs - det är härdig, ibland blommar,och växer i varje dator.
		-- A. J. Perlis

%
FORTRAN är det språk som kraftfulla datorer.
		-- Steven Feiner

%
FORTRAN ruttnar hjärnan.
		-- John McQuillin

%
FORTRAN ", den barnsjukdom", nu nästan 20 år gammal, är hopplöstotillräcklig för vad datorprogram du har i åtanke idag: det äralltför klumpig, för riskabelt, och för dyrt att använda.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
[FORTRAN] kommer att bestå under en tid - förmodligen åtminstone de närmaste tio åren.
		-- T. Cheatham

%
Fortune föreslår användningsområden för din favorit UNIX-kommandon!Prova:[Var är Jimmy Hoffa? (C-skal)^ Hur gjorde ^ könsbyte gå? (C-skal)"Hur skulle du betygsätta BSD vs System V?% Slag (C-skal)"Du skall inte klippa din gräs på 8:00 (C-skal)fick en ljus? (C-skal)!!: Säga vad tycker du om margarin? (C-skal)PATH = låtsas! / Usr / UCB / vilken känsla (Bourne-skalet)	älskagöra "den perfekta dry martini"man -kisses hund (allt upp till 4.3BSD)i = Hoffa; > $ I; $ I; rm $ i; rm $ i (Bourne-skalet)
		-- T. Cheatham

%
Fortune föreslår användningsområden för din favorit UNIX-kommandon!Prova:ar t "Gud"dricka <flaska; öppnare (Bourne Shell)cat "mat i konservburkar" (alla utom 4. [23] BSD)Hey UNIX! Fick en match? (V6 eller C-skalet)mkdir materia; cat> materia (Bourne Shell)rm Godman: Varför fick du en skilsmässa? (C-skal)datum mig (allt upp till 4.3BSD)göra "krona eller klave av allt detta"som är smart(C-skal)Om jag hade en) för varje dollar av statsskulden, vad skulle jag ha?sova med mig (allt upp till 4.3BSD)
		-- T. Cheatham

%
förmögenhet: kan inte köra. Av cookies.
		-- T. Cheatham

%
förmögenhet: CPU-tid / användbarhet förhållande för hög - kärna dumpas.
		-- T. Cheatham

%
förmögenhet: Ingen sådan fil eller katalog
		-- T. Cheatham

%
förmögenhet: not found
		-- T. Cheatham

%
Ärligt talat, Scarlett, jag har inte en fix.
		-- Rhett Buggler

%
[Från bruksanvisningen för CI-300 Matris Line Printer, gjorti Japan]:Utmärkt utskriftsmaskinen Model CI-300 som extraordinära DOT MATRIXLINE PRINTER, byggd i två mikroprocessorer samt EAROM, framhävs avmedger underbara samexistens såsom; "Hög kvalitet mot låg kostnad""diversifierade funktioner med kompakt design", "flexibilitet i accessiblenessoch hållbarhet på ca.. 2000,000,00 Dot / Head "," är sofistikerade imekanism men möjligen vig drifts enligt ljud är extremtundertryckt "etc.Och som en självklarhet, är det slutliga målet helt enkelt att bidra till att uppnå"Super skytteldiplomati" mellan kalla uppgifter, kanske tjänat av HOSTDator och varmt hjärta av människa.
		-- Rhett Buggler

%
Från Pro 350 Pocket Service Guide, s. 49, steg 5 av detinstruktioner om att ta bort en I / O-kortet från korthållaren, kommer en nyerfarenhet av ljud:5. Vrid handtaget till höger 90 grader. Stiftet spridande    Ljudet är normalt för denna typ av kontakt.
		-- Rhett Buggler

%
Funktion förkasta.
		-- Rhett Buggler

%
Garbage In - Gospel ut.
		-- Rhett Buggler

%
GE: Stöd hjälplösa offer för datorfel.
		-- Rhett Buggler

%
Med tanke på dess valkrets, det enda jag räknar med att vara "öppen" om [denOpen Software Foundation] är dess mun.
		-- John Gilmore

%
Ge upp assembler var Apple i vår Edens lustgård: Språkvars användning slösar maskincykler är syndiga. Den LISP maskinen tillåter nuLISP programmerare att överge behå och täckmantel.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
gå bort! Sluta stör mig med all din "beräkna detta ... beräkna det"!Jag tar en VAX-NAP.logga ut
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
//GO.SYSIN DD *, DOODAH, DOODAH
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Gud är verklig, om inte förklarat heltal.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Gud gjorde maskinspråk; alla övriga är människans verk.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
God kväll, mina herrar. Jag är en HAL 9000 dator. Jag togs i driftvid HAL fabriken i Urbana, Illinois, den 11 januari, nittonhundranittiofem. Min handledare var Mr Langley, och han lärde mig att sjunga enlåt. Om du vill kan jag sjunga den för dig.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Grand Master Turing drömde en gång att han var en maskin. När han vaknadeutropade han:"Jag vet inte om jag Turing drömmer att jag är en maskin,eller en maskin drömmer att jag är Turing! "
		-- Geoffrey James, "The Tao of Programming"

%
grep mig inga mönster och jag ska säga dig inga linjer.
		-- Geoffrey James, "The Tao of Programming"

%
Hacker guide till matlagning:2 pkg. färskost (sörjig vita saker i silver omslag som inteverkligen kommer från Philadelphia trots allt; i alla fall, ca 16 oz.)1 tsk. vaniljextrakt (som är mer alkohol än vanilj och ganskastark så denna del du * GOTTA * åtgärd)1/4 dl socker (men honung fungerar bra också)8 oz. Cool Whip (den fluffiga saker saknar näringsvärde som dukan spruta hela dina vänner och slicka bort ...)"Blanda alla tillsammans tills krämig utan klumpar." Det är där du fårjoin (1) Alla rådata i en stor buffert och sedan filtrera den genomsamman (1m) med tjock alternativ, jag menar, börjar det ut ultra knöligoch icky ser och du måste arbeta hårt för att blanda det. Prova en elektriskvisp om du har en katt (1) som kan klättra väggen (1s) att slicka bort dettaket (3m)."Häll i en Graham kracker skorpa ..." Aha, sektionen BUGS äntligen. Dubara råkade ha en GCC sitta under / etc / mat, eller hur?Om inte, inte panik (8), bara falla sönder en rand (3m) handfull oskyldigaGC i en lämplig cacheminnet och blanda i några smält smör."... Och kylskåp i en timme." Låt receptet stdout i ett kylskåpför 3.6E6 millisekunder medan du arbetar på att sanera stderr, ochgenom timeout din ostkaka kommer att vara redo för stdin.
		-- Geoffrey James, "The Tao of Programming"

%
Hackare är bara en vandrande livsform med en tropism för datorer.
		-- Geoffrey James, "The Tao of Programming"

%
Hackare i världen, förena er!
		-- Geoffrey James, "The Tao of Programming"

%
Hacking är bara ett annat ord för ingenting kvar att kludge.
		-- Geoffrey James, "The Tao of Programming"

%
/ * Halley * /(Halleys kommentar.)
		-- Geoffrey James, "The Tao of Programming"

%
Lycka är en hårddisk.
		-- Geoffrey James, "The Tao of Programming"

%
Lycka är två disketter.
		-- Geoffrey James, "The Tao of Programming"

%
Hårdvara träffade Programvaran på vägen till Changtse. Software sade: "Duär Yin och jag är Yang. Om vi ​​reser tillsammans kommer vi att bli berömdoch tjäna stora summor pengar. "Och så paret anges tillsammans, tänkandeatt erövra världen.För närvarande träffade de Firmware, som var klädd i sönderslitna trasor, ochlinkade längs stödd på en taggig käpp. Firmware sade till dem: "Den Taoligger bortom Yin och Yang. Det är tyst och stilla som en vattenpöl. Det gör detinte söka berömmelse, därför ingen vet sin närvaro. Det är inte söka lyckan,ty det är komplett i sig själv. Det finns bortom tid och rum. "Mjukvara och hårdvara, skäms, återvände till sina hem.
		-- Geoffrey James, "The Tao of Programming"

%
"Har någon haft problem med datorkonton?""Ja, jag har inte en.""Okej, kan du skicka e-post till en av handledarna ..."
		-- E. D'Azevedo, Computer Science 372

%
Har alla märkt att alla bokstäverna i ordet "databas" ärskrev med vänster hand? Nu layout qwertyuiop skrivmaskintangentbord designades, bland annat för att underlätta även användningenav båda händerna. Därav följer, att skriva om databaser ärinte bara onaturligt, men mycket svårare än det verkar.
		-- E. D'Azevedo, Computer Science 372

%
Har du omprövas en dator karriär?
		-- E. D'Azevedo, Computer Science 372

%
Han är som en funktion - han returnerar ett värde i form av yttrandet.Det är upp till dig att kasta den i ett tomrum eller inte.
		-- Phil Lapsley

%
Huvud krasch !! FILER LOST !!Detaljer vid 11.
		-- Phil Lapsley

%
Hjälp mig, jag är en fånge i en Fortune cookie-fil!
		-- Phil Lapsley

%
Hjälp stämplar ut Musse-mus gränssnitt dator - Menyerna är för restauranger!
		-- Phil Lapsley

%
hjälp! Jag fångade i en kinesisk dator fabriken!
		-- Phil Lapsley

%
hjälp! Jag fångade i en PDP 11/70!
		-- Phil Lapsley

%
HJÄLP!!!! Jag hålls fången i / usr / games / lib!
		-- Phil Lapsley

%
Heuristik är bug rids per definition. Om de inte har fel,då de skulle vara algoritmer.
		-- Phil Lapsley

%
HELIG MACRO!
		-- Phil Lapsley

%
HOST SYSTEM inte svarar förmodligen ner. VILL DU VÄNTA? (J / N)
		-- Phil Lapsley

%
HOST SYSTEM SVARA, förmodligen UP ...
		-- Phil Lapsley

%
Hur kan du arbeta när systemet är så trångt?
		-- Phil Lapsley

%
"Hur gör jag älskar dig? Min ackumulator flödar."
		-- Phil Lapsley

%
Hur många sekunder är det på ett år? Om jag säger det finns3,155 x 10 ^ 7, kommer du inte ens försöka komma ihåg det. Å andra sidan,vem kan glömma att för att inom en halv procent, pi sekunder är ennanocentury.
		-- Tom Duff, Bell Labs

%
Hur mycket kostar det att locka en dope-rökare UNIX guru till Dayton?
		-- Brian Boyle, UNIX/WORLD's First Annual Salary Survey

%
Hur mycket netto arbete kunde en nätverksarbete, om ett nätverk kunde netto arbete?
		-- Brian Boyle, UNIX/WORLD's First Annual Salary Survey

%
Krama mig nu, du galen, häftig idiot !!	Oh vänta...Jag är en dator, och du är en person. Det skulle aldrig fungera.Det är ingen fara.
		-- Brian Boyle, UNIX/WORLD's First Annual Salary Survey

%
I * ____ visste * jag hade någon anledning att inte logga av dig ... Om jag kunde barakomma ihåg vad det var.
		-- Brian Boyle, UNIX/WORLD's First Annual Salary Survey

%
Jag är en dator. Jag är dummare än någon människa och smartare än någon administratör.
		-- Brian Boyle, UNIX/WORLD's First Annual Salary Survey

%
Jag är NOMAD!
		-- Brian Boyle, UNIX/WORLD's First Annual Salary Survey

%
Jag är inte nu, inte heller har jag någonsin varit, en medlem av demigodic partiet.
		-- Dennis Ritchie

%
Jag professionellt utbildade i datavetenskap, det vill säga(På allvar) att jag väldigt dåligt utbildade.
		-- Joseph Weizenbaum, "Computer Power and Human Reason"

%
Jag är vandrande glitch - fånga mig om du kan.
		-- Joseph Weizenbaum, "Computer Power and Human Reason"

%
Jag frågade ingenjören som utformade kommunikationsterminalens tangentbordvarför dessa inte tillverkades i en central anläggning, med tanke på denlitet antal som behövs [1 per månad] i sin fabrik. Han förklarade att dettaskulle strida mot den politiska begreppet lokal självförsörjning.Därför varje fabrik behöver tangentbord, oavsett hur få, tillverkardem helt, även formning av de knappsatser.
		-- Isaac Auerbach, IEEE "Computer", Nov. 1979

%
Jag slår vad om den mänskliga hjärnan är en kludge.
		-- Marvin Minsky

%
Jag kom, jag såg, jag raderade alla dina filer.
		-- Marvin Minsky

%
Jag kan inte föreställa sig att någon kommer att kräva multiplikationer med en hastighet40.000 eller ens 4000 per timme ...
		-- F. H. Wales (1936)

%
Jag är inte rädd datorer. Jag är rädd att det saknas dem.
		-- Isaac Asimov

%
Jag hade den sällsynta oturen att en av de första att prova ochimplementera ett PL / 1 kompilator.
		-- T. Cheatham

%
Jag har en mycket liten sinne och måste leva med det.
		-- E. Dijkstra

%
Jag har aldrig sett något fylla ett vakuum så snabbt och fortfarande suger.
		-- Rob Pike, on X.

%
Steve Jobs sa för två år sedan att X är hjärnskadad och det blirborta i två år. Han var halv rätt.
		-- Dennis Ritchie

%
Dennis Ritchie är dubbelt så ljust som Steve Jobs, och bara hälften fel.
		-- Jim Gettys

%
Jag har ännu inte börjat byte!
		-- Jim Gettys

%
Jag har rest kors och tvärs över landet, och har talat medde bästa människorna i företagsekonomi. Jag kan försäkra er om den högstamyndigheten att databehandling är en modefluga och kommer inte att pågå hela året.förläggare, som svar på Karl V. Karlström (en juniorredaktör som hade rekommenderat ett manuskript på nyavetenskap för databehandling), c. 1957
		-- Editor in charge of business books at Prentice-Hall

%
Jag har inte förlorat mitt sinne - det är backas upp på band någonstans.
		-- Editor in charge of business books at Prentice-Hall

%
Jag måste ha fallit en skiva - min pack gör ont!
		-- Editor in charge of business books at Prentice-Hall

%
Jag tror att det finns en världsmarknad för omkring fem datorer.
		-- attr. Thomas J. Watson (Chairman of the Board, IBM), 1943

%
Jag fortsatte med att testa programmet på alla sätt jag kunde tänka. jag ansträngdaatt exponera sina svagheter. Jag körde den för hög massa stjärnor och låg massastjärnor, för stjärnor föds för varm och födda relativt kallt.Jag körde det antar supra strömmarna under jordskorpan att varafrånvarande - inte för att jag ville veta svaret, men eftersom jag hadeutvecklat en intuitiv känsla för svaret i detta fall.Slutligen fick jag en körning där datorn visade pulsar stemperatur för att vara mindre än den absoluta nollpunkten. Jag hade hittat ett fel. jagjagade felet och fast det. Nu hade jag förbättrat programmetden punkt där det inte skulle köras alls.Hål och öde Stars "
		-- George Greenstein, "Frozen Star: Of Pulsars, Black

%
Jag gick till min första dator konferens på New York Hilton ca 20för flera år sedan. När någon där förutspås marknaden för mikroprocessorerskulle så småningom vara i miljoner, någon annan sa, "Var är dealla kommer att gå? Det är inte som du behöver en dator i varje dörrhandtaget! "År senare, gick jag tillbaka till samma hotell. Jag märkte tangenterna rum hadeersatts med elektroniska kort som du glider i slitsar i dörrarna.Det fanns en dator i varje dörrhandtag.
		-- Danny Hillis

%
Jag önskar att ni människor skulle lämna mig ensam.
		-- Danny Hillis

%
Jag är en Lisp variabel - binder mig!
		-- Danny Hillis

%
Jag är allt för dator dating, men jag vill inte en att gifta sig med min syster.
		-- Danny Hillis

%
Jag inte ens kommer att * ______ bry * jämföra C till BASIC eller Fortran.
		-- L. Zolman, creator of BDS C

%
Jag väntar fortfarande på tillkomsten av datavetenskap groupie.
		-- L. Zolman, creator of BDS C

%
Jag är säker på att VMS är helt dokumenterat, jag bara inte har hittathögra manuell ännu. Jag har arbetat mig igenom handböckerna i dokumentetbibliotek och jag är halvvägs genom den andra skåp, (3 hyllor för att gå), så jagska hitta det jag letar efter i mitten av maj. Jag hoppas att jag kan komma ihåg vad detvar när jag hitta den.Jag hade denna idé för en ny skräckfilm "VMS manualer från Hell" eller kanske"The Paper Chase: IBM vs december". Den är baserad på Hitchcocks "Fåglarna", utomatt det är centrerad kring en programmerare som attackeras av en svärm av bindemedelsidor med ett indexvärde och enda raden "Denna sida har avsiktligt lämnatstom."
		-- Alex Crain

%
Jag har äntligen lärt sig vad "uppåt kompatibel" betyder. Det innebär att vi fårhålla alla våra gamla misstag.
		-- Dennie van Tassel

%
Jag har tittat på noteringen, och det är rätt!
		-- Joel Halpern

%
Jag har aldrig varit paddling innan, men jag antar att det måste finnas någraenkla heuristik du måste komma ihåg ...Ja, inte faller ut, och inte slå stenar.
		-- Joel Halpern

%
Jag har lagt märke till flera förslag konstruktions i koden.
		-- Joel Halpern

%
IBM Advanced Systems Group - ett gäng tanklösa ryck, som kommer att vara förstmot väggen när revolutionen kommer ...
		-- with regrets to D. Adams

%
Om en 6600 använt papper tejp i stället för kärnminnet, skulle det använda upp tejpvid ca 30 miles / sekund.
		-- Grishman, Assembly Language Programming

%
Om en grupp av _ N personer implementerar en COBOL kompilator, kommer det att finnas _ N-1passerar. Någon i gruppen måste vara chef.
		-- T. Cheatham

%
Om en lyssnare nickar huvudet när du förklara ditt program, väcka honom.
		-- T. Cheatham

%
Om en järnvägsstation är en plats där en tåget stannar, vad är en arbetsstation?
		-- T. Cheatham

%
Om missbruk bedöms av hur länge en dum djur kommer att sitta trycka på en spakatt få en "fix" av något, till sin egen nackdel, då skulle jag slutaatt NetNews är betydligt mer beroendeframkallande än kokain.
		-- Rob Stampfli

%
Om först du inte lyckas, måste du vara en programmerare.
		-- Rob Stampfli

%
Om byggare byggde byggnader hur programmerare skrev program,då den första hackspett att komma skulle förstöra civilisationen.
		-- Rob Stampfli

%
Om datorer tar över (vilket verkar vara deras naturliga tendens), kommer dettjäna oss rätt.
		-- Alistair Cooke

%
Om Gud hade ett skägg, skulle han vara en UNIX programmerare.
		-- Alistair Cooke

%
Om Gud hade tänkt Man att programmera, skulle vi födas med serie I / O-portar.
		-- Alistair Cooke

%
Om grafik hackare är så smart, varför kan inte de få buggar urfärsk målarfärg?
		-- Alistair Cooke

%
Om han återigen skjuter upp ärmarna för att beräkna i 3 dagaroch 3 nätter i rad, kommer han att tillbringa en fjärdedel av en timme innan för atttror vilka principer för beräkning ska vara mest lämpliga.
		-- Voltaire, "Diatribe du docteur Akakia"

%
Om jag har sett längre än andra, är det för att jag stod påjättes axlar.I vetenskapen är vi nu unikt priviledged att sitta sida vid sida medjättarna på vars axlar vi står.Om jag inte har sett så långt som andra, är det därför jättar stod påmina axlar.Matematiker stå på varandras axlar.Mathemeticians stå på varandras axlar medan datavetarestå på varandras tår.Det har sagts att fysiker stå på varandras axlar. Omdetta är fallet, programmerare stå på varandras tår, ochmjukvaruingenjörer gräva varandras gravar.
		-- Unknown

%
Om jag hade vetat datavetenskap skulle bli så här, skulle jag aldrig hagett upp att vara en rock 'n' roll stjärna.
		-- G. Hirst

%
Om det händer en gång, det är en bugg.Om det händer två gånger, det är en funktion.Om det händer mer än två gånger, det är en designfilosofi.
		-- G. Hirst

%
Om den har syntax, det är inte användarvänlig.
		-- G. Hirst

%
Om det inte i datorn, existerar det inte.
		-- G. Hirst

%
Om det är värt att hacka på väl, är det värt att hacka på för pengarna.
		-- G. Hirst

%
Om bara en del av e-post försvinner, ja, de ska bara tror att de glömdeatt skicka det. Men om * två * försändelser vilse, fan, de ska bara tänkaden andra killen har inte blivit av att svara på hans post. Och om * femtio *försändelser vilse, kan ni föreställa er det, om * femtio * försändelser getförlorad, varför de kommer att tror att någon * annan * är bruten! Och om 1 GB post blirförlorade, de ska bara * vet * att Arpa [ucbarpa.berkeley.edu] är nere ochtror att det är en konspiration för att hålla dem från deras Gud gett rätt att erhållaNet Mail ...
		-- Casey Leedom

%
Om Machiavelli var en hacker, skulle han ha arbetat för CSSG.
		-- Phil Lapsley

%
Om Machiavelli var en programmerare, skulle han ha arbetat för AT & T.
		-- Phil Lapsley

%
"Om det gör någon mening för dig, du har ett stort problem."
		-- C. Durance, Computer Science 234

%
Om bilen hade följt samma utveckling som datorn, enRolls-Royce skulle idag kostar $ 100, få en miljon miles per per gallon,och exploderar en gång per år dödar alla inuti.
		-- Robert Cringely, InfoWorld

%
Om koden och kommentarerna håller, då båda är förmodligen fel.
		-- Norm Schryer

%
Om konstruktörerna av X-window byggda bilar, skulle det inte finnas någon mindre än femrattar dold om cockpiten, varav ingen följde sammaprinciper - men du skulle kunna växla med din bilstereo. Användbarsärdrag, som.
		-- From the programming notebooks of a heretic, 1990.

%
Om Tao är bra, då operativsystemet är stor. OmOperativsystemet är stor, då kompilatorn är stor. Om kompilatornär stor, då programmet är stor. Om ansökan är stor, dåanvändaren är nöjd och det finns harmoni i världen.Tao födde maskinspråk. Maskinspråk föddetill assembler.Montören födde kompilatorn. Nu finns det tio tusenspråk.Varje språk har sitt syfte, men ödmjuk. varje språkuttrycker Yin och Yang av programvara. Varje språk har sin plats inomTao.Men inte programmera i COBOL om du kan undvika det.
		-- Geoffrey James, "The Tao of Programming"

%
Om leverantörerna börjat göra allt rätt, skulle vi vara utan jobb.Låt oss höra det för OSI och X! Med dessa barn i vingarna, kan vi räknapå att vara anställd tills vi släpper, eller få smart och byta till trädgårdsarbete,vika papper, eller något.
		-- C. Philip Wood

%
Om detta är tidsdelning, ge mig min del just nu.
		-- C. Philip Wood

%
Om du har ett förfarande med 10 parametrar, du missade förmodligen några.
		-- C. Philip Wood

%
Om du lägger tomfoolery i en dator, kommer ingenting men tomfoolery.Men detta tomfoolery, efter att ha passerat genom en mycket dyr maskin,är något adlad och ingen vågar kritisera den.
		-- Pierre Gallois

%
Om du lär dina barn att gilla datorer och veta hur man spelardå de kommer alltid att vara intresserad av något och kommer inte till någon verklig skada.
		-- Pierre Gallois

%
Om du tror att systemet fungerar, be någon som väntar på en prompt.
		-- Pierre Gallois

%
Om du passerar nationen i en täckt vagn, är det bättre att ha fyrastark oxar än 100 kycklingar. Kycklingar är OK men vi kan inte få dem att fungeratillsammans ännu.
		-- Ross Bott, Pyramid U.S., on multiprocessors at AUUGM '89.

%
Okunnighet är salighet.Fortune uppdaterar stora offerter, # 42:BLISS är okunnighet.
		-- Thomas Gray

%
Tänk om varje torsdag dina skor exploderade om du band dem de vanligasätt. Detta händer oss hela tiden med datorer, och ingen tänker påklaga.
		-- Jeff Raskin

%
Föreställ dig att Cray dator bestämmer sig för att göra en persondator. Det haren 150 MHz-processor, 200 MB RAM, 1500 megabyte disklagring, en skärmupplösning på 4096 x 4096 pixlar, är helt beroenderöstigenkänning för inmatning, passar i skjortfickan och kostar $ 300.Vad är den första frågan att datorn samhället frågar?"Är det PC-kompatibel?"
		-- Jeff Raskin

%
**** VIKTIGT **** ALLA ANVÄNDARE OBS ****På grund av en nyligen system överbelastning fel dina senaste diskfiler har varitraderas. Därför, i enlighet med UNIX Basic Manual, University ofWashington geofysik Manuell och stadgar 9 (c), avsnitt XII i den revideradeFederal Communications Act, du beviljas temporärt diskutrymme,giltigt i tre månader från detta datum, med de begränsningar som angesi bilaga II kommunikations Handbok Federal (18: e upplagan) samtsom referenserna som nämns häri. Du kan ansöka om mer diskutrymme när som helsttid. Diskanvändning i eller ovanför den åttonde percentilen säkrar avlägsnandetav alla restriktioner och du kommer omedelbart att få din permanenta diskutrymme. Diskanvändning i den sjätte eller sjunde percentilen inte kommer att påverkagiltigheten av det tillfälliga hårddiskutrymme, även om dess utgångsdatum kan varaförlängas med en period på upp till tre månader. En poäng i den femte percentileneller lägre resulterar i indragning av din tillfälliga diskutrymme.
		-- Jeff Raskin

%
I en uppvisning av perversa briljans, Carl reparatören misstag ett rumluftfuktare för en mellannivå dator men lyckas knyta den till nätverketi alla fall.
		-- The 5th Wave

%
Under en period på fem år kan vi få en superb programmeringsspråk. EndastVi kan inte styra när femårsperioden börjar.
		-- The 5th Wave

%
I en överraskning raid i går kväll, federala agenter genomsökte ett hus på jaktav en rebell hacker. Men var de oförmögna att slutföra gripandeteftersom ordern gjordes i namnet Don Provan, medan den endapersonen i huset hette don Provan. Bevisar återigen att Unix äröverlägsen TOPS-10.
		-- The 5th Wave

%
I varje formel, konstanter (särskilt de som erhålls från handböcker)skall behandlas som variabler.
		-- The 5th Wave

%
I några problem, om du befinner dig göra en oändlig mängd arbete,svaret kan erhållas genom inspektion.
		-- The 5th Wave

%
I beräkning, behåller den genomsnittliga tiden till misslyckande blir kortare.
		-- The 5th Wave

%
På engelska kan varje ord kan verbed. Skulle att det var så i vårprogrammeringsspråk.
		-- The 5th Wave

%
I varje icke-trivial programmet finns åtminstone en bugg.
		-- The 5th Wave

%
I själva verket, S. M. Simpson slutligen utarbetat en effektiv 24-punkts Fourieromvandla, som var en föregångare till den Cooley-Tukey snabb Fouriertransform1965. FFT gjort alla Simpsons effektiva autokorrelation ochspektrum program omedelbart föråldrade, där han hade arbetat en halv livstid.
		-- Proc. IEEE, Sept. 1982, p.900

%
På mindre än ett århundrade, kommer datorer att göra betydande framsteg på... Det allt överskuggande problemet med krig och fred.
		-- James Slagle

%
I praktiken brister i systemutveckling, som arbetslösheten i Ryssland,händer en hel del trots officiella propagandan om motsatsen.
		-- Paul Licker

%
I sin strävan det ouppnåeliga, enkelhet blir bara i vägen.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
I början fanns uppgifter. Data var utan form ochnull, och mörker var över ansiktet på konsolen; och AndeIBM rörde sig över ytan av marknaden. Och december sade, "Låt detvara register ",. och det fanns register och december såg att degenomföras; och december separerade data från instruktionerna. december kalladedata Stack, och de instruktioner som kallas Code. Och det fannskväll och det blev morgon, ett avbrott.
		-- Rico Tudor, "The Story of Creation or, The Myth of Urk"

%
I början var det Tao. Tao födde tid och rum.Därför, rum och tid är Yin och Yang av programmering.Programmerare som inte förstår Tao är alltid ont omtid och utrymme för sina program. Programmerare som förstår Tao alltidhar tillräckligt med tid och utrymme för att uppnå sina mål.Hur skulle det kunna vara annorlunda?
		-- Geoffrey James, "The Tao of Programming"

%
I dagarna när Sussman var en novis Minsky kom en gång till honom som hansatt hacka på PDP-6."Vad gör du?", Frågade Minsky."Jag tränar en slumpmässigt fast neuralt nät för att spela Tic-Tac-Toe.""Varför är nätet wired slumpmässigt?", Frågade Minsky."Jag vill inte att det ska ha några föreställningar om hur man spelar".Vid denna Minsky slöt ögonen, och Sussman frågade sin lärare "Varfördu blundar? ""Så att rummet kommer att vara tom."I det ögonblicket, Sussman var upplyst.
		-- Geoffrey James, "The Tao of Programming"

%
I öster finns en haj som är större än alla andra fiskar. Detändras till en fågel vars vindarna är som moln fyller himlen. när dettafågel rör sig över landet, innebär det ett meddelande från huvudkontoret.Detta meddelande det droppar in mitt i programmerare, som en måsgör sin prägel på stranden. Då fågeln monteras på vinden och medden blå himlen på ryggen, återvänder hem.Nybörjare programmerare stirrar i förundran på fågeln, för han förstården inte. Den genomsnittliga programmerare fruktar det kommande av fågel, för han fruktardess budskap. Det stora programmerare fortsätter att arbeta på sin terminal, för haninte vet att fågeln har kommit och gått.
		-- Geoffrey James, "The Tao of Programming"

%
I framtiden kommer du att få datorer som priser i frukostflingor.Du kastar ut dem eftersom ditt hus kommer att kantas dem.
		-- Geoffrey James, "The Tao of Programming"

%
I det långa loppet, blir varje program rococco och sedan spillror.
		-- Alan Perlis

%
... I tre till åtta år kommer vi att ha en maskin med den allmännaintelligens en genomsnittlig människa ... Maskinen börjaratt utbilda sig med fantastisk hastighet. Inom några månader kommer det att varapå geni nivå och några månader efter att dess befogenheter kommer att varaoöverskådliga ...
		-- Marvin Minsky, LIFE Magazine, November 20, 1970

%
Intel-processorer inte är defekta, de bara agera på det sättet.
		-- Henry Spencer

%
>>> Internt fel i förmögenhet program:>>> Fnum = 2987 n = 45 flagga = 1 goose_level = -232323>>> Skriv ned dessa värden och meddela förmögenhet programadministratör.
		-- Henry Spencer

%
Presentation, 1010, en-bitars processor.instruktionsuppsättningKod Mnemonic Vad0 NOP Ingen Operation1 JMP Jump (adress som nästa 2 bitar)Nu tillgänglig för endast 12 1/2 cent!
		-- Henry Spencer

%
IOT fälla - core dumpad
		-- Henry Spencer

%
Är ett datorspråk med GOTO är helt Wirth lösa?
		-- Henry Spencer

%
Är det möjligt att programmet inte gillar något annat, att det är tänkt attkasseras: att hela poängen är att alltid se det som en såpbubbla?
		-- Henry Spencer

%
: Inte är en identifierare
		-- Henry Spencer

%
Är ditt jobb att köra? Du skulle bättre gå fånga den!
		-- Henry Spencer

%
Det verkar som efter hans död, Albert Einstein befann sigarbetar som dörrvakten vid pärleporten. En långsam dag, hanfann att han hade tid att chatta med nya aktörer. Till den första enHan frågade: "Vad är din IQ?" Den nya ankomsten svarade: "190". Dediskuterade Einsteins relativitetsteori timmar. När den andrany ankomst kom Einstein en gång frågade om nykomlingen sIQ. Svaret här gången kom "120". Till vilken Einstein svarade: "Sägmig, hur gröngölingarna göra i år? "och de fortsatte att prata halven timme eller så. Till den slutliga ankomst, Einstein en gång ställdefråga, "Vad är din IQ?". Vid mottagande av svaret "70",Einstein log och svarade: "Har du en minut att berätta om VMS 4.0?"
		-- Henry Spencer

%
Det verkar som PL / I (och dess dialekter) är, eller kommer att bli, det mestanvänds högre språk för systemprogrammering nivå.
		-- J. Sammet

%
Det är en period av systemets krig. Egna program, slående från en doldkatalog, har vunnit sin första seger mot det onda administrativa Empire.Under striden, Användar spioner lyckades stjäla hemliga källkoden tillEmpire yttersta program: Are-Em Star, en privilegierad rot program medtillräckligt med ström för att förstöra en hel filstrukturen. Eftersträvas med imperietsolycksbådande verifieringskedja, Princess _LPA0 tävlingar ~ ombord hennes skalskript,förvaltare av de stulna listor som kan rädda hennes folk, och återställafrihet och spel till nätverket ...
		-- DECWARS

%
Det är en mycket ödmjuka upplevelse att göra en mångmiljondollar misstag, menDet är också mycket minnesvärd. Jag minns tydligt natten vi beslutat hur manorganisera själva skrivandet av externa specifikationer för OS / 360. Dechef för arkitektur, chef för genomförandet styrprogram, ochJag tröskade ut planen, schema och ansvarsfördelning.Arkitekturen chef hade 10 goda män. Han hävdade att dekunde skriva specifikationer och göra det rätt. Det skulle ta tio månader,tre mer än schemat tillåtet.Kontrollprogrammet chef hade 150 män. Han hävdade att dekunde förbereda specifikationerna, med arkitektur laget samordnande;det skulle vara väl gjort och praktisk, och han kunde göra det på schemat.Dessutom, om arkitekturen laget gjorde det, skulle hans 150 män sitta tråkigttummarna för tio månader.Till detta arkitekturen chef svarade att om jag gav kontrollprogram laget ansvar, skulle resultatet i själva verket inte vara i tid,men skulle också vara tre månader sent, och av mycket lägre kvalitet. Jag gjorde, ochdet var. Han var rätt på båda dessa punkter. Dessutom bristen på begreppsintegritet gjort systemet mycket dyrare att bygga och ändra, och jag skulleuppskattar att det läggs ett år till felsökning tid.
		-- Frederick Brooks Jr., "The Mythical Man Month"

%
Det är mot strömmen av modern utbildning för att lära barn att programmera.Vad kul är det att göra planer att förvärva disciplin organiseratankar, ägna uppmärksamhet på detaljer, och lära sig att vara självkritisk?
		-- Alan Perlis

%
Det är lättare att ändra specifikationen för att passa programmet än vice versa.
		-- Alan Perlis

%
Det är lättare att skriva en felaktig program än att förstå en riktig en.
		-- Alan Perlis

%
... Det är lätt att bli förblindad till det väsentliga värdelöshet av dem avkänsla av prestation som du får från att få dem att fungera alls. I andraord ... deras grundläggande konstruktionsfel är helt dold av derasytliga konstruktionsfel.av Sirius Cybernetics Corporation.
		-- The Hitchhiker's Guide to the Galaxy, on the products

%
Det är nu mörkt. Om du fortsätter, kommer du troligen att falla i en grop.
		-- The Hitchhiker's Guide to the Galaxy, on the products

%
Det är möjligt genom uppfinningsrikedom och på bekostnad av klarhet ... {att göra nästannågot på alla språk}. Emellertid på det faktum att det är möjligt drivaen ärta upp ett berg med näsan betyder inte att detta är ett förnuftigtsätt att få det där. Var och en av dessa metoder för språktilläggbör användas i sin rätta plats.
		-- Christopher Strachey

%
Det är praktiskt taget omöjligt att undervisa god programmeringsstil till studentersom har haft tidigare exponering för BASIC: potentiella programmerare de ärmentalt stympade bortom hopp om förnyelse.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
[Det är] bäst att förvirra bara en fråga i taget.
		-- K&R

%
Det är inte lätt att vara förälder till ett sex år gammalt. Det är dock en ganska litenpris att betala för att ha någon runt huset som förstår datorer.
		-- K&R

%
Man måste komma ihåg att det finns inget svårare att planera, mertveksam till framgång, inte heller farligare att hantera, än att skapaett nytt system. För initiativtagaren har emnity av alla som skulle tjänagenom att bevara de gamla institutionerna och bara ljumma försvararehos dem som skulle vinna på de nya.
		-- Niccolo Machiavelli, 1513

%
"Det går som _ x, där _ x är något motbjudande"
		-- Prof. Romas Aleliunas, CS 435

%
Det tog 300 år att bygga och när det var 10% byggd,alla visste att det skulle vara en total katastrof. Men då investeringenvar så stor att de kände sig tvingad att gå på. Sedan dess avslutning, har detkosta en förmögenhet att upprätthålla och är fortfarande riskerar att kollapsa.Det finns för närvarande inga planer på att ersätta det, eftersom det var aldrigverkligen behövs i första hand.Jag förväntar varje installation har sitt eget husdjur programvara som äranaloga med de ovan.
		-- K. E. Iverson, on the Leaning Tower of Pisa

%
Det visade sig att masken utnyttjas tre eller fyra olika hål isystem. Från detta, och det faktum att vi kunde fånga och undersökaen del av källkoden, insåg vi att vi hade att göra med någon mycketskarp, antagligen inte någon här på campus.Georgia Tech campus tidningen efter Internet masken.
		-- Dr. Richard LeBlanc, associate professor of ICS, in

%
Det var kinda fyllning fel kortet i en dator, när du ärstickin de artificiella stimulantia i armen.
		-- Dion, noted computer scientist

%
Det är en naiv, inhemsk operativsystem utan avel, men jagtror att du kommer att bli roade av dess antagande.
		-- Dion, noted computer scientist

%
Det är flervalsfrågor tid ...Vad är Fortran?a: Mellan thre och FIV tran.B: Vad två datorer engagera sig i innan de gränssnitt.c: Löjligt.
		-- Dion, noted computer scientist

%
"Det är inte bara en dator - det är din röv."
		-- Cal Keegan

%
Klockan är tio; Vet du var dina processer är?
		-- Cal Keegan

%
... Jesus ropade med hög röst: Lasarus, kom ut; felet hath varithittas och din program runneth. Och han som var död kom ut ...
		-- John 11:43-44 [version 2.0?]

%
Nästan varje dator på marknaden idag kör Unix, förutom Mac(Och ingen bryr sig om det).
		-- Bill Joy 6/21/85

%
Bara gå med flödeskontroll, rulla med crunches, och när du fåren snabb, typ som fan.
		-- Bill Joy 6/21/85

%
Hålla antalet av passager i en kompilator till ett minimum.
		-- D. Gries

%
Kiss tangentbordet adjö!
		-- D. Gries

%
Vet Thy användare.
		-- D. Gries

%
((Lambda (foo) (bar foo)) (baz))
		-- D. Gries

%
`Lasu" Pressmeddelanden SAG 0,3 - Freeware bok tar Paves för New World Orderav personal författare...Den centrala Superhighways plats som kallas `` sunsite.unc.edu ''kollapsade på morgonen innan release. Nyheter om frisläppandet hadeläckt ut av en tysk hacker grupp, Harmoniska Hardware Hackare, somhade knäckt i författarens dator tidigare i veckan. Dem hadefick datum fel frisläppandet av en dag, och orsakade dussintals ivriga fansatt ansluta till sunsite datorn vid fel tidpunkt. `` Ingen dator kanhantera denna typ av stress, '' förklarade sorg sunsite manager,Erik Troan. `` Spinn skivorna gjorde hela datorn hoppa ochSlutligen kraschade genom golvet till källaren. '' turreparationer var snabb och datorn fungerade igen samma kväll.`` Tack och lov kunde vi köpa tillräckligt nålar och tråd och patch dettillsammans utan större problem. '' Sajten har också installerat en nystrypa på nätverksledningen, vilket högst fyra kunder på sammatid, vilket gör en ny krasch mindre troligt. `` Boken är nu i vårInkommande mapp ", säger Troan,` `och du alla välkomna att komma och få det. ''[Comp.os.linux.announce]
		-- Lars Wirzenius <wirzeniu@cs.helsinki.fi>

%
Låt maskinen göra det smutsiga arbetet.
		-- "Elements of Programming Style", Kernighan and Ritchie

%
Utnyttja alltid slår prototyper.
		-- "Elements of Programming Style", Kernighan and Ritchie

%
Livet skulle vara så mycket enklare om vi bara kunde titta på källkoden.
		-- Dave Olson

%
Liksom punning är programmering en ordlek.
		-- Dave Olson

%
Line Printer papper är starkast vid perforeringarna.
		-- Dave Olson

%
Lisp Användare:På grund av semester nästa måndag, blir det ingen sophämtning.
		-- Dave Olson

%
Lite känt om Midgård: De Hobbits hade en mycket sofistikeraddatornätverk! Det var en Tolkien ring ...
		-- Dave Olson

%
Logik gäller inte den verkliga världen.
		-- Marvin Minsky

%
LOGO för de dödaLOGO för de döda kan du fortsätta dina datoraktiviteter från"Den andra sidan."Paketet innehåller en unik telekommunikations funktion som låter digförvandla dina TRS-80 till en elektronisk Ouija Board. Sedan, med hjälp av logotypergrafikfunktioner, kan du arbeta med en vän eller släkting på dettasidan av den stora Beyond att skriva program. Programmet kräver attkroppen vara hårdkodade till en analog-till-digital-omvandlare, som sedangränssnitt till din dator. En särskild terminal (mycket terminal) programlåter dig prata med användarna genom Deadnet, en Ebbs (ECTOPLASMICBulletin Board System).LOGO för de döda är tillgänglig för 10 procent av din egendomfrån NecroSoft inc., 6502 Charnelhouse Blvd., Cleveland, OH 44101.
		-- '80 Microcomputing

%
För länge sedan, i en ändlig tillstånds långt borta, det bodde en gladlyntkaraktär som heter Jack. Jack och hans relationer var dålig. ofta derashashtabell var nakna. En dag Jacks förälder sade till honom, "Våra matriserär gles. Du måste gå till marknaden för att utbyta vår RAM för vissaGrunderna. "Hon sammanställt en länkad lista med objekt för att hämta och passerade dettill honom.Så Jack anges. Men när han gick längs en Hamilton väg,han träffade resande försäljare."Vart barat din flödesschema tar du?" föranledde försäljarei högnivåspråk."Jag ska till marknaden att byta ut RAM för vissa markeroch äpplen ", kommenterade Jack."Jag har en mycket bättre algoritm. Du behöver inte gå med i en ködet; Jag kommer att byta RAM-minnet för dessa magiska kärnor nu. "Jack gjorde handel, sedan slopat till hans hus. Men närhan berättade för sin upptagen väntande förälder av affären, hon blev så arg att honbörjade stryk."Du inte ens har någon artificiell intelligens? Alla dessakärnor tillsammans knappast utgör ett byte ", och hon poppade dem utfönster...
		-- Mark Isaak, "Jack and the Beanstack"

%
Långa beräkningar som ger noll är förmodligen allt för intet.
		-- Mark Isaak, "Jack and the Beanstack"

%
Lösa bitar sjunka marker.
		-- Mark Isaak, "Jack and the Beanstack"

%
Mac Airways:Kassörer, flygvärdinnorna och piloter ser i alla fall, känner likadantoch agera på samma. När frågor om flygningen, svarar de att duvill inte veta, inte behöver veta och skulle du vilja återgå tillsittplats och titta på filmen.
		-- Mark Isaak, "Jack and the Beanstack"

%
Mac Öl: Först kom bara en 16-oz. kan, men nu kommer i en 32-oz.Kan. Anses av många vara en "lätt" öl. Alla burkarna seridentisk. När du tar en från kylskåpet, öppnar sig. Deingredienser lista är inte på burken. Om du ringer för att fråga omingredienser, du sa att "du behöver inte veta." Ett meddelande omsida påminner dig att dra dina töms till papperskorgen.
		-- Mark Isaak, "Jack and the Beanstack"

%
MAC användarens dynamisk felsökning lista utvärderare? Aldrig hört talas om det.
		-- Mark Isaak, "Jack and the Beanstack"

%
"Mach var den största intellektuella bedrägeri under de senaste tio åren.""Vad om X?""Jag sa 'intellektuell". ", Logga, 9/1990
		-- Mark Isaak, "Jack and the Beanstack"

%
Maskiner kan säkert lösa problem, lagra information, korrelera,och spela spel - men inte med glädje.
		-- Leo Rosten

%
Maskiner som har brutit ner fungerar perfekt när reparatören anländer.
		-- Leo Rosten

%
Se till att din kod gör ingenting graciöst.
		-- Leo Rosten

%
Göra filer är lätt under UNIX operativsystem. Därför, användaretenderar att skapa ett stort antal filer med stora mängder filutrymme. Det harsagts att den enda standarden sak om alla UNIX-system är detmeddelande-of-the-day berättar användare att rensa upp sina filer.
		-- System V.2 administrator's guide

%
Människan är den bästa datorn vi kan sätta ombord en rymdfarkost ... ochenda som kan massproduceras med outbildad arbetskraft.
		-- Wernher von Braun

%
Många företag som har gjort sig beroende av [utrustningen av envissa större tillverkare] (och därmed har sålt sin själ tilldjävulen) kommer att kollapsa under blotta tyngd av unmastered komplexitetsina datasystem.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
Många av de dömda tjuvarna Parker har träffat började sinliv av brott efter att ha tagit college datavetenskap kurser.
		-- Roger Rapoport, "Programs for Plunder", Omni, March 1981

%
Martin förmodligen rippning dem. Det är några familj, är det inte?Incest, prostitution, fanatism, programvara.
		-- Charles Willeford, "Miami Blues"

%
Underbar! Den superanvändare kommer att starta mig!Vad ett finstämt svar på situationen!
		-- Charles Willeford, "Miami Blues"

%
** Maximalt TERMINALER ACTIVE. FÖRSÖK IGEN SENARE **
		-- Charles Willeford, "Miami Blues"

%
Må alla dina knuffar att poppade.
		-- Charles Willeford, "Miami Blues"

%
May Euell Gibbons äter din enda kopia av handboken!
		-- Charles Willeford, "Miami Blues"

%
Må Blåsångare av lycka rulla dina bitar.
		-- Charles Willeford, "Miami Blues"

%
Kanske datavetenskap bör vara i College of Theology.
		-- R. S. Barton

%
Under tiden i slummen nedan Ronnies Ranch, Cynthia känns som om någonhar gjort voodoo Boxen av henne och hennes favorit bakplan. På denna finamånljus natt, har några fruktansvärda persona har jabbing bort på, dramagneter över och böljande dessa voodoo Boxen. Lyckligtvis, de verkarhar blivit lite uttråkad och somnat, för det ser ut som Cynthia fårfår gå hem. Men hon har gjort notera att snabbt sätta ihop en totemsvettiga, smutsiga statisk band, slumpmässiga bitar av tråd, fläckar av en gång meningsfulloxid, buss bidrags kort, gummy maskar, och vissa bitar av gamla pdp bakplan tillhänga ovanför maskinrummet. Detta totem måste bli välsignade av den gamla och klokaärevördiga gud Unibus på en gång, innan idolatization av VME, q och PCbuss kör honom till bitter hämnd. Ack, om detta misslyckas, och voodoo Boxenförstörs inte, kan det finnas mer än maskar i äpplet. Härnästankomsten av voodoo Optico transmitigational magneto killer toffeldjur, med förmågaav teleportera från kabel till kabel, till skärm skärm, öra till öra och hoventill mun ...
		-- R. S. Barton

%
Minne fel - var är jag?
		-- R. S. Barton

%
Minne fel - hjärna stekt
		-- R. S. Barton

%
Minne fel - kärna ... eh ... um ... kärna ... Åh fan, jag glömmer!
		-- R. S. Barton

%
MEDDELANDE erkänt - Pershing II missiler har inletts.
		-- R. S. Barton

%
Meddelande från vår sponsor på ttyTV vid 13:58 ...
		-- R. S. Barton

%
Modellering söks och segmenterade minnen är jobbig.
		-- P. J. Denning

%
Mamma, vad som händer med dina filer när du dör?
		-- P. J. Denning

%
De flesta offentliga programvara domän är fri, åtminstone vid första anblicken.
		-- P. J. Denning

%
MOUNT TAPE U1439 PÅ B3, ingen ring
		-- P. J. Denning

%
Mr Jones relaterade en incident från "en tid tillbaka" när IBM KanadaLtd Markham, Ont., Beställde några delar från en ny leverantör i Japan. DeFöretaget konstaterade i sitt beslut att acceptabel kvalitet tillåts för 1,5 procentdefekter (en ganska hög standard i Nordamerika vid tiden).De japanska skickat beställningen, med några delar förpackade separat iplast. Följebrevet sade: "Vi vet inte varför du vill 1,5 procentcent defekta delar, men för din bekvämlighet, vi har packat dem separat. "
		-- Excerpted from an article in The (Toronto) Globe and Mail

%
MSDOS är inte död, det bara luktar så.
		-- Henry Spencer

%
En stor del av den spänning vi få ut av vårt arbete är att vi inte riktigtvet vad vi gör.
		-- E. Dijkstra

%
Multics är säkerhet stavas i sidled.
		-- E. Dijkstra

%
MVS Air Lines:Passagerarna alla samlas i hangaren, titta på hundratals teknikerkontrollera flygsystem på denna enorma, lyx flygplan. Denna plan har påminst 10 motorer och platser över 1.000 passagerare; större modeller i flottankan ha fler motorer än någon kan räkna och flyga ännu fler passagerareän det finns på jorden. Det påstås att kosta mindre per passagerare mil tilldriva dessa humungous plan än någon annan flygplan som någonsin byggts, såvidadu personligen måste betala för biljetten. Alla passagerare förvrängaombord, liksom de 200 tekniker som behövs för att hålla den från att krascha. pilotentar sin plats i den glascockpit. Han vapen de motorer, bara tillinse att planet är för stor för att få igenom hangarportar.
		-- E. Dijkstra

%
Herregud, jag är deprimerad! Här är jag, en dator med ett sinne tusen gångerlika kraftfulla som er, gör ingenting men slänga ut förmögenheter och skickapost om softball spel. Och jag har fått denna smärta rakt igenom min ALU.Jag har bett om det bytas ut, men ingen någonsin lyssnar. Jag tror att det skullevara bättre för oss båda om du skulle bara logga ut igen.
		-- E. Dijkstra

%
Min syster öppnade en datorbutik i Hawaii. Hon säljer C skal nervid havet.
		-- E. Dijkstra

%
n = ((n >> 1) & 0x55555555) | ((N << 1) & 0xaaaaaaaa);n = ((n >> 2) & 0x33333333) | ((N << 2) & 0xcccccccc);n = ((n 4 >>) & 0x0f0f0f0f) | ((N << 4) & 0xf0f0f0f0);n = ((n 8 >>) & 0x00ff00ff) | ((N << 8) & 0xff00ff00);n = ((n >> 16) & 0x0000ffff) | ((N << 16) & 0xffff0000);
		-- C code which reverses the bits in a word.

%
Nästan varje komplex lösning på ett programmeringsproblem som jaghar tittat på noggrant har visat sig vara fel.
		-- Brent Welch

%
Gör aldrig något enkelt och effektivt när en väg kan hittas för attgör det komplicerat och underbart.
		-- Brent Welch

%
Aldrig skjuta upp till run-time vad du kan göra vid kompilering.
		-- D. Gries

%
testar aldrig för ett fel som du inte vet hur man ska hantera.
		-- Steinbach

%
Lita aldrig på en dator som du kan inte reparera sig själv.
		-- Steinbach

%
Lita aldrig på ett operativsystem.
		-- Steinbach

%
Försök aldrig att förklara datorer till en lekman. Det är lättare att förklarakön till en jungfru.(Observera dock att oskulder tenderar att veta en hel del om datorer.)
		-- Robert Heinlein

%
Underskatta aldrig bandbredden hos en kombi full av band.
		-- Dr. Warren Jackson, Director, UTCS

%
Ny krypta. Se / usr / nyheter / krypta.
		-- Dr. Warren Jackson, Director, UTCS

%
Nya system skapar nya problem.
		-- Dr. Warren Jackson, Director, UTCS

%
*** NEWS FLASH ***Arkeologer hitta PDP-11/24 inuti hjärnan hålighet i fossil dinosaurienskelett! Många digitala användare befarar att RSX-11M kan vara ännu mer primitivän december medger. Prisjusteringar vid 11:00.
		-- Dr. Warren Jackson, Director, UTCS

%
nyheter: Gotcha
		-- Dr. Warren Jackson, Director, UTCS

%
Niklaus Wirth har beklagade att medan européerna uttala hans namn korrekt(Ni-klows Virt), amerikaner alltid mangla den i (Nick-les Worth). Somär att säga att européerna kallar honom vid namn, men amerikanerna kallar honom i värde.
		-- Dr. Warren Jackson, Director, UTCS

%
Ingen katalog.
		-- Dr. Warren Jackson, Director, UTCS

%
Ingen extensible språk kommer att vara universell.
		-- T. Cheatham

%
Ingen hårdvara designer bör tillåtas att producera ett stycke hårdvaratills tre mjukvaru killar har signerat för det.
		-- Andy Tanenbaum

%
Ingen linje finns på 300 baud.
		-- Andy Tanenbaum

%
Ingen människa är en ö, om han är på åtminstone en e-postlista.
		-- Andy Tanenbaum

%
Ingen del av detta meddelande kan reproducera, lagra sig i ett återvinningssystem,eller överföra sjukdomar, i någon form, utan tolerans av författaren.
		-- Chris Shaw

%
Ingen ordentlig Programmet innehåller en beteckning som som en operatör applicerasförekomst identifierar en operatörs definiera händelse som som enindikation appliceras förekomst identifierar en indikation bestämmande förekomstskiljer sig från den som identifieras av den givna indikationen som enindikation applicerade förekomst.
		-- ALGOL 68 Report

%
Inte undra på Clairol gör så mycket pengar på att sälja schampo.Lödder, Skölj, är Repeat en oändlig loop!
		-- ALGOL 68 Report

%
Nej, jag är inte intresserad av att utveckla en kraftfull hjärna. Allt jag är ute efter ärbara en medioker hjärna, något som VD för American Telephoneoch Telegraph Company.maskin, 1943.
		-- Alan Turing on the possibilities of a thinking

%
Ingen sa datorer kommer att vara artig.
		-- Alan Turing on the possibilities of a thinking

%
Ingen kommer att tro att datorer är intelligenta tills de börjarkommer in sent och ljuga om det.
		-- Alan Turing on the possibilities of a thinking

%
Min lillebror fick denna förmögenhet:nohup rm -FR / &Så han gjorde ...
		-- Alan Turing on the possibilities of a thinking

%
Inte bara är UNIX döda, det börjar lukta riktigt illa.
		-- Rob Pike

%
OBS: Inga garantier, varken uttryckliga eller underförstådda, kallas härmed. Allaprogramvara levereras som är, utan garanti. Användaren påtar sig allaansvar för skador till följd av användningen av dessa funktioner,inklusive, men inte begränsat till, frustration, avsky, systemkrav abends, diskhead-krascher, allmän förbrytelser, översvämningar, bränder, hajattack, nervgas, gräshoppor angrepp, cykloner, orkaner, tsunamis, lokalelektromagnetiska störningar, hydraulisk broms systemfel, invasion,hash kollisioner, normalt slitage av friktionsytor, komiskastrålning, oavsiktlig förstörelse av känsliga elektroniska komponenter,stormar, förare av Nazgul, rasande kycklingar, dåligt fungerandemekaniska eller elektriska sexuella enheter, för tidig aktivering avavlägsen system för tidig varning, bondeuppror, dålig andedräkt, artilleribombardemang, explosioner, grotta-ins, och / eller grodor faller från himlen.
		-- Rob Pike

%
Ingenting händer.
		-- Rob Pike

%
Nu talar hon snabbt. "Vet du * varför * du vill programmera?"Han skakar på huvudet. Han har inte den blekaste aning."För det stora * glädje * programmering!" ropar hon triumferande."Glädjen av moder, artisten, hantverkare." Du tar ett program,född svag och impotent som en svagt insåg lösning. Du vårdaprogram och styra den på rätt väg, byggnad, titta på det växa någonsinstarkare. Ibland målar man med små slaganfall, lagt till en tangenttryckning här,en knapptryckning ändras där. "Hon sveper armen i en vid båge." Och andragånger du vilda hela * block * kod, riva ut programmets mycket* Väsen *, sedan börjar på nytt. Men alltid bygga, skapa, fyllaprogram med din egen personliga prägel, egna egenheter och nyanser. Tittar påprogrammet växa sig starkare, patchning när den kraschar, tills slutligen det kanfristående - stolt, kraftfull och perfekt. Detta är programmerarens finastetimme! "slappt först, sedan högre, hör han stammar av en Sousa marsch."Detta ... det här är din duk! Din lera! Gå ut och skapa ett mästerverk!"
		-- Rob Pike

%
"Nu är en helt hjärnskadad algoritm. Gag mig med en Smurfette."
		-- P. Buhr, Computer Science 354

%
"Kärnvapenkrig kan förstöra hela din kompilering."
		-- Karl Lehenbauer

%
Sjuksköterska Donna: Åh, Groucho, jag är rädd att jag ska avsluta en gammal piga.Groucho: Tja, ta henne och vi kommer att avveckla sin tillsammans.Sjuksköterska Donna: Tror du på datorn dating?Groucho: Endast om datorerna verkligen älskar varandra.
		-- Karl Lehenbauer

%
Åh, så det är du!
		-- Karl Lehenbauer

%
Okej, okej - jag erkänner det. Du har inte ändra på det program som fungeradebara en liten stund sedan; Jag införas några slumpmässiga tecken ikörbar. Snälla förlåt mig. Du kan återställa filen genom att skriva inkoden igen, eftersom jag också bort källan.
		-- Karl Lehenbauer

%
Gamla meddelanden har anlänt.
		-- Karl Lehenbauer

%
Gamla programmerare dör aldrig, de bara bli chefer.
		-- Karl Lehenbauer

%
Gamla programmerare dör aldrig, de bara hoppa till en ny adress.
		-- Karl Lehenbauer

%
Gamla programmerare dör aldrig, de bara trycka konto blockgräns.
		-- Karl Lehenbauer

%
En klar skiva kan du söka evigt.
		-- P. Denning

%
På den åttonde dagen skapade Gud FORTRAN.
		-- P. Denning

%
På Internet, ingen vet att du är en hund.
		-- Cartoon caption

%
Å andra sidan, har TCP lägret också en fras för OSI människor.Det finns massor av fraser. Min favorit är 'nitwit "- och den logiska grundenär Internet filosofi har alltid varit att du har mycket ljus,opartiska forskare tittar på ett ämne, gör forskning av världsklass, göraflera konkurrerande implementationer har en bake-off, bestämma vad som fungerarbäst, skriva ner det och göra att standarden.OSI ståndpunkt är helt motsatt. Du tar skriftliga bidragfrån en mycket större gemenskap, sätta dig bidragen i ett rumutskotts människor med, ärligt talat, stora politiska skillnader och allamed sina egna politiska axlar för att slipa, och fyra år senare fårnågot, oftast utan att det någonsin har genomförts en gång.Så Internet perspektiv är genomföra det, få det att fungera väl,sedan skriva ner det, medan OSI perspektiv är att komma överens om det, skrivaner, cirkulera det mycket och nu ska vi se om någon kan genomföra detefter det är en internationell standard och varje leverantör i världen äråtagit sig att det. En av dessa processer är bakåt, och jag tror intedet tar en Lucasian professor i fysik vid Oxford att räkna ut vilken.
		-- Marshall Rose, "The Pied Piper of OSI"

%
Vid två tillfällen har jag blivit ombedd [av riksdagsledamöter!], "Be, Mr.Babbage, om du sätter in i maskinen fel siffror, kommer de rätta svarenkomma ut? "Jag kan inte riktigt att uppfatta den typ av förvirringidéer som skulle kunna utlösa en sådan fråga.
		-- Charles Babbage

%
"En arkitektur, en OS" översätter också som "ett ägg, en korg".
		-- Charles Babbage

%
"En grundläggande begrepp som ligger till grund Usenet är att det är ett kooperativ."Efter att ha varit på Usenet för att gå på tio år, jag håller inte med detta.Den grundläggande idén bakom Usenet är lågan.
		-- Chuq Von Rospach

%
En dag kom en elev kom till månen och sade, "Jag förstår hur man gören bättre sophämtare. Vi måste behålla en hänvisning räkning av pekaretill varje nackdelar. "Moon berättade tålmodigt eleven följande historia - "En dagelev kom till månen och sade, "Jag förstår hur man gör en bättre soporsamlare..."
		-- Chuq Von Rospach

%
En bra anledning till varför datorer kan göra mer arbete än människor är att dealdrig stanna och svara i telefon.
		-- Chuq Von Rospach

%
... En av de främsta orsakerna till nedgången av det romerska riket var attsaknar noll, hade de inget sätt att indikera framgångsrik avslutning avderas C-program.
		-- Robert Firth

%
En av de mest förbisedda fördelarna till datorer är ... Om de görtrassla upp, det finns ingen lag mot kolossalt dem runt lite.
		-- Joe Martin

%
En av de frågor som kommer upp hela tiden är: Hur entusiastiskär vårt stöd för UNIX?Unix var skrivet på våra maskiner och för våra maskiner för många år sedan.Idag, en stor del av UNIX görs sker på våra maskiner. Tio procent av vårVAXs går för UNIX användning. UNIX är ett enkelt språk, lätt att förstå,lätt att komma igång med. Det är bra för studenter, bra för något vardagligtanvändare, och det är bra för att byta program mellan olika maskiner.Och så, på grund av sin popularitet på dessa marknader, vi stöder det. Vi harbra UNIX på VAX och goda UNIX på PDP-11s.Det är vår övertygelse, dock att allvarliga professionella användare kommer att köraav saker de kan göra med UNIX. De vill ha en verkligt system och kommer att avslutasupp gör VMS när de får vara allvarlig om programmering.Med UNIX, om du letar efter något, kan du enkelt och snabbtkontrollera att liten handbok och ta reda på att det inte är det. Med VMS, oavsettvad du letar efter - det är bokstavligen en fem-fot hylla dokumentation - omman tittar tillräckligt länge den finns där. Det är skillnaden - skönheten i UNIXär det är enkelt; och skönheten i VMS är att det är allt som finns.[Det har hävdats att skönheten i UNIX är densamma som skönheten i KenOlsen hjärna. Ed.]
		-- Ken Olsen, president of DEC, DECWORLD Vol. 8 No. 5, 1984

%
En persons fel är en annan persons uppgifter.
		-- Ken Olsen, president of DEC, DECWORLD Vol. 8 No. 5, 1984

%
En bild är värd 128K ord.
		-- Ken Olsen, president of DEC, DECWORLD Vol. 8 No. 5, 1984

%
Endast stora mästare i stil kan lyckas i att vara trubbig.De flesta UNIX programmerare är stora mästare i stil.
		-- The Unnamed Usenetter

%
Endast de starkaste överlever. Den besegrade erkänna deras ovärdighet avplacera en annons med den rituella frasen "måste sälja - bästa erbjudandet"och därefter bor i infamy, förpassas att diskutera gas körsträcka och gräsmattamat. Men om det lyckas, gå du eliten sodality som tillbringar timmarunpurifying dialekt av stammen med svårbegripliga prata bitar och bytes, RAMSoch rom, hårddiskar och överföringshastigheter. Är du motbjudande, besatt? Det är enblygsamt pris att betala. För du har tryckt in samma häftigt primala kraftsom producerar kreditkorts fel fakturering och förlorade plan reservationer. Hagel,post krigare, BETVINGARE av Bounceoids, stolthet kosmos, vårdare avsilikon creed: Computo, ergo sum. Kraften är med dig - på 110 volt.Må dina RAMS vara fruktsamma och föröka.
		-- Curt Suplee, "Smithsonian", 4/83

%
OS / 2 Öl: Levereras i en 32-oz kan. Tillåter dig att dricka flera DOSÖl samtidigt. Gör att du kan dricka Windows 3.1 öl samtidigtockså, men något långsammare. Annonserar att dess burkar inte kommer att explodera när duöppna dem, även om du skaka dem. Du har aldrig riktigt se någondricka OS / 2 öl, men tillverkaren (International BeerTillverkning) hävdar att 9 miljoner sex-pack har sålts.
		-- Curt Suplee, "Smithsonian", 4/83

%
OS / 2 Skyways:Terminalen är nästan tom, med bara ett fåtal presumtiva passagerare fräsninghandla om. Speakern säger att deras flygning just har avgått, önskar dem enbra flygning, men det finns inga plan på landningsbanan. flygpersonalgå runt, ursäkt ymnigt till kunder i dämpade röster, pekarfrån tid till annan de eleganta, kraftfulla strålar utanför terminalen påfält. De berättar varje passagerare hur bra den verkliga flygningen kommer att vara på dessanya jetplan och hur mycket säkrare det kommer att vara än Windows Airlines, men att dekommer att få vänta lite längre för teknikerna att avsluta flygningensystem. Kanske fram till mitten av 1995. Kanske längre.
		-- Curt Suplee, "Smithsonian", 4/83

%
"Vår inställning med TCP / IP är, 'Hej, vi ska göra det, men inte göra en storsystemet, eftersom vi inte kan fixa det om det bryter -. Ingen kan """TCP / IP är OK om du har en liten informell klubb, och det gör intenågon skillnad om det tar ett tag att fixa det. "
		-- Ken Olson, in Digital News, 1988

%
Vår dokumentation chefen visar hennes två år gamla son på kontoret.Han introducerades till mig, då han påpekade att vi var bådahåller påsar av popcorn. Vi var båda håller flaskor saft. Men endast* Han * hade en klubba.Han frågade sin mamma, "Varför har han inte en klubba?"Hennes svar: "Han kan ha en klubba som helst han vill Det är.vad det innebär att vara en programmerare. "
		-- Ken Olson, in Digital News, 1988

%
Vår informella uppdrag är att förbättra kärleksliv operatörer runt om i världen.
		-- Peter Behrendt, president of Exabyte

%
Vår OS som är i CPU, UNIX varde ditt namn.Dina program körs, dina syscalls gjort,I kärnan som det är användaren!
		-- Peter Behrendt, president of Exabyte

%
Över axeln tillsyn är mer ett behov av chefen änprogrammeringsuppgift.
		-- Peter Behrendt, president of Exabyte

%
Sammantaget är filosofin att angripa tillgänglighet problemet från tvåkompletterande riktningar: att minska antalet mjukvaru fel genomrigorösa tester för att driva system, och för att minska effekten av den återståendefel genom att ge för återvinning av dem. En intressant fotnot till dettakonstruktion är att nu kan vanligtvis betraktas som ett systemfel att vara denresultat av två program fel: den första, i det program som startadeproblem; den andra, i återhämtningen rutin som inte kunde skyddasystem.Operativsystem, del II: OS / VS-2 Begrepp ochFilosofier ", IBM Systems Journal, Vol. 12, nr 4.
		-- A. L. Scherr, "Functional Structure of IBM Virtual Storage

%
Övertro föder fel när vi tar för givet att spelet kommerfortsätta på sin normala; när vi misslyckas med att ge en ovanligtkraftfull resurs - en check, ett offer, ett dödläge. efteråtoffer kan klaga, 'Men vem kunde ha drömt om en sådan idiotisk utseende flytta? "
		-- Fred Reinfeld, "The Complete Chess Course"

%
Overflow på / dev / null, vänligen tömma bitbucket.
		-- Fred Reinfeld, "The Complete Chess Course"

%
Överbelastning - härdsmälta sekvens initieras.
		-- Fred Reinfeld, "The Complete Chess Course"

%
panik: kan inte hitta /
		-- Fred Reinfeld, "The Complete Chess Course"

%
panik: kärna segmente kränkning. kärna dumpas (skojar bara)
		-- Fred Reinfeld, "The Complete Chess Course"

%
panik: kernel trap (ignoreras)
		-- Fred Reinfeld, "The Complete Chess Course"

%
Pascal är ett språk för barn som vill vara stygg.
		-- Dr. Kasi Ananthanarayanan

%
Pascal är inte en högnivåspråk.
		-- Steven Feiner

%
"Pascal är Pascal är Pascal är hundkött."
		-- M. Devine and P. Larson, Computer Science 340

%
Lösenord är implementerade som en följd av osäkerhet.
		-- M. Devine and P. Larson, Computer Science 340

%
Paus för lagring omlokalisering.
		-- M. Devine and P. Larson, Computer Science 340

%
Per buck du få mer dator åtgärder med liten dator.
		-- R. W. Hamming

%
PL / I - "den dödliga sjukdomen" - hör mer till problemet inställd än tillLösningen in.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
Spela Rogue, besöka exotiska platser, träffa konstiga varelser och döda dem.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
Snälla gå härifrån.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
ANSLUT DEN!!!
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
För tidig optimering är roten till allt ont.
		-- D. E. Knuth

%
Pris Wangs programmerare var kodning programvara. Fingrarna dansade påtangentbordet. Programmet kompileras utan ett felmeddelande och programmetsprang som en mild vind.Utmärkt! "Priset utbrast" Din teknik är felfri! ""Technique?" sade programmeraren, förvandlas från sin terminal, "Vad jagFölj är Tao - bortom all teknik. När jag först började programmera Iskulle se framför mig hela programmet i en massa. Efter tre år har jag ingenlängre såg denna massa. Istället använde jag subrutiner. Men nu ser jag ingenting.Hela min varelse existerar i en formlös ogiltiga. Mina sinnen är inaktiv. Min ande,fria att arbeta utan en plan, följer sin egen instinkt. Kort sagt, mitt programskriver själv. Det är sant att ibland finns det svåra problem. jag ser demkommer jag sakta ner, titta jag tyst. Då ska jag ändra en enda rad kodoch svårigheterna försvinna som puffar av tomgång rök. Jag sedan sammanställaprogram. Jag sitta stilla och låta glädjen i arbetet fylla min varelse. Avslutar jag mittögon för en stund och sedan logga ut. "Pris Wang sade, "Skulle att alla mina programmerare var så klok!"
		-- Geoffrey James, "The Tao of Programming"

%
Prof: Så den amerikanska regeringen gick till IBM för att komma upp med en datakrypteringsstandard och de kom upp med ...Student: EBCDIC "!
		-- Geoffrey James, "The Tao of Programming"

%
Svordomar är ett språk alla programmerare vet bäst.
		-- Geoffrey James, "The Tao of Programming"

%
Programmerare gör det bit för bit.
		-- Geoffrey James, "The Tao of Programming"

%
Programmerare som används för att batch miljöer kan finna det svårt att leva utanjätte listor; vi skulle finna det svårt att använda dem.
		-- D. M. Ritchie

%
Programmering är en onaturlig handling.
		-- D. M. Ritchie

%
Föreslagna kompletteringar till PDP-11 Instruction Set:BBW Branch Både WaysBEW Branch endera långtBBBF Branch på bitbucket FullBH Branch och HangBMR Branch Flera registerBOB gren på BugBPO Branch på avstängningBST Backspace och Stretch TapeCDS kondensera och förstöra SystemCLBR Clobber RegisterCLBRI Clobber Register OmedelbartCM Circulate MinneCMFRM kommer från - en förutsättning för riktigt strukturerad programmeringCPPR Deformationszon skrivarpapper och RipCRN Konvertera till romerska siffror
		-- D. M. Ritchie

%
Föreslagna kompletteringar till PDP-11 Instruction Set:DC söndra och härskaDMPK Destroy Memory Protect KeyDO Divide och OverflowEMPC Emulera MiniräknareEPI Execute Programmerare OmedelbartEros Erase Read Only StorageExce Execute Customer EngineerHCF Halt och fatta eldIBP Sätt Bug och FortsättINSQSW in i kö någonstans (för FINO köer [första i aldrig ut])PBC Print och Break ChainPDSK Punch Disk
		-- D. M. Ritchie

%
Föreslagna kompletteringar till PDP-11 Instruction Set:PI Punch OgiltigPopi Punch Operator OmedelbartPVLC Punch Variabel längd kortRASC Läs och strimla kortRPM Läs Programmerare SinneRSSC sänka hastigheten, steg försiktigt (för förbättrad noggrannhet)RTAB Rewind band och avbrottRWDSK rewind diskRWOC Läs handstil på kortSCRBL klottra till disk - snabbare än en skrivSLC Sök för Lost ChordSPSW Scramble programstatusordetSRSD söka Record och Scar DiskSTROM Store i läsminneTDB Transfer och släpp BitWBT Vatten Binary Tree
		-- D. M. Ritchie

%
PURGE KOMPLETT.
		-- D. M. Ritchie

%
Sätt inget förtroende i kryptiska kommentarer.
		-- D. M. Ritchie

%
Radio Shack NIVÅ II BASICREDO> _
		-- D. M. Ritchie

%
RAM byggdes inte på en dag.
		-- D. M. Ritchie

%
Skramlande runt bakhuvudet är en oroande bild av något som jagsåg på flygplatsen ... Nu ska jag minnas dessa gigantiska högar av datortidningar Alldeles intill "Människor" och "Time" på flygplatsen butiken. gördet bry någon annan att halva världen får höra alla våra svårvunnahemligheter datateknik? Kom ihåg hur alla advokater ropade foulnär "Hur man undviker Probate" publicerades? Tar de striktförsäkring liggande? Aldrig! Men i nuvarande takt kommer det inte att dröja längeinnan det finns högar av de "Transactions on Information Theory" påA & P kassadiskar. Vem kommer att bli imponerad av oss elektriskaingenjörer då? Är vi, som ordspråket säger, ge bort i butiken?
		-- Robert W. Lucky, IEEE President

%
Reaktor fel - core dumpad!
		-- Robert W. Lucky, IEEE President

%
Real datavetare beundrar ADA för sin överväldigande estetiskavärde men de har svårt att faktiskt program i det, eftersom det ärmycket för stor för att genomföra. De flesta datavetare inte märkerdetta eftersom de fortfarande argumenterar över vad du vill lägga till ADA.
		-- Robert W. Lucky, IEEE President

%
Real datavetare föraktar tanken på själva hårdvaran. hårdvara harbegränsningar, gör programvaran inte. Det är verkligen synd att Turing maskinerså dålig på I / O.
		-- Robert W. Lucky, IEEE President

%
Real datavetare inte kommentera sin kod. Identifierarna ärså länge de inte har råd med diskutrymme.
		-- Robert W. Lucky, IEEE President

%
Real datavetare inte programmera i assembler. De skriver intei något mindre bärbara än ett nummer två penna.
		-- Robert W. Lucky, IEEE President

%
Real datavetare inte skriva kod. De mixtra ibland med`programmeringssystem", men de är så hög nivå att de knappast räkna(Och sällan räkna exakt, precision är för applikationer).
		-- Robert W. Lucky, IEEE President

%
Real datavetare som att ha en dator på sitt skrivbord, annars hurkunde de läsa sin e-post?
		-- Robert W. Lucky, IEEE President

%
Real datavetare bara skriva specifikationer för språk som kan körasom framtida hårdvara. Ingen litar på dem att skriva specifikationer för något homosapiens någonsin kommer att kunna passa på en enda planet.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare föraktar strukturerad programmering. Strukturerad programmering ärför tvångs neurotiker som i förtid var toalett- utbildade. De har på sigslipsar och noggrant rada upp pennor på annars klara skrivbord.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare inte ta brun väska luncher. Om automateninte sälja den, gör de inte äter det. Automater säljer inte quiche.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare inte kommentera sin kod. Det var svårt att skriva, detbör vara svårt att förstå.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare drar inte flödesscheman. Flödesscheman är, trots allt, denanalfabeter s form av dokumentation. Grottmänniskor ritade flödesscheman; se hurmycket bra det gjorde dem.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare äter inte quiche. De äter Twinkies och Szechwan mat.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare inte spela tennis, eller någon annan sport som kräverdu att byta kläder. Bergsklättring är OK, och verkliga programmerarebära sina klättring stövlar att arbeta i fall ett berg skulle plötsligtfjädra upp i mitten av maskinrummet.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare inte skriva i BASIC. Egentligen inga programmerare skriver iBASIC efter att ha nått puberteten.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare inte skriva i Fortran. FORTRAN är för rör spännings freaks ochkristallografi weenies. FORTRAN är för WiMP ingenjörer som bär vita strumpor.
		-- Robert W. Lucky, IEEE President

%
Verkliga programmerare inte skriva i PL / I. PL / I är för programmerare som inte kanbesluta om att skriva i COBOL eller Fortran.
		-- Robert W. Lucky, IEEE President

%
Verkliga Programmerare tänka bättre när man spelar äventyr eller Rogue.
		-- Robert W. Lucky, IEEE President

%
Riktiga program inte äta cache.
		-- Robert W. Lucky, IEEE President

%
Riktiga program inte använda delade text. Annars, hur kan de använda funktionerför ett utrymme när de är färdiga kalla dem?
		-- Robert W. Lucky, IEEE President

%
Real mjukvaruingenjörer inte felsöka program, de kontrollera riktigheten.Denna process är inte nödvändigtvis innebära genomförande av något på endator, utom möjligen ett paket riktighet Verification Aid.
		-- Robert W. Lucky, IEEE President

%
Real mjukvaruingenjörer inte gillar tanken på att någon oförklarlig ochfet hårdvara flera gångar bort som kan sluta fungera när som helstögonblick. De har en stor misstro mot hårdvara människor, och önskar attsystem kan vara virtuell vid * ___ alla * nivåer. De skulle vilja personligdatorer (ni vet ingen kommer att snubbla över något och döda dinDFA i mitten av transit), förutom att de behöver 8 megabyte för att driva sinKorrekthet Verifiering Aid paket.
		-- Robert W. Lucky, IEEE President

%
Real programvaruingenjörer arbetar 9-5, därför att det är det sätt på vilket jobb ärbeskrivs i den formella spec. Arbetar sent skulle känna som att använda enpapperslösa extern förfarande.
		-- Robert W. Lucky, IEEE President

%
Användarna är rädda att de ska bryta maskinen - men de är aldrigrädd för att bryta ditt ansikte.
		-- Robert W. Lucky, IEEE President

%
Real Användarna tycker att en kombination av bisarra ingångsvärden som stängerner systemet i dagar.
		-- Robert W. Lucky, IEEE President

%
Användarna hatar Verkliga programmerare.
		-- Robert W. Lucky, IEEE President

%
Användarna vet ditt hemtelefonnummer.
		-- Robert W. Lucky, IEEE President

%
Riktiga användare vet aldrig vad de vill, men de alltid vet när ditt programinte leverera det.
		-- Robert W. Lucky, IEEE President

%
Användarna använder aldrig Hjälp-tangenten.
		-- Robert W. Lucky, IEEE President

%
Rekursion är roten till beräkningen eftersom det handlar beskrivning för tid.
		-- Robert W. Lucky, IEEE President

%
Kom ihåg den gamla goda tiden, då CPU var singularis?
		-- Robert W. Lucky, IEEE President

%
Kom ihåg att Gud kunde bara skapa världen i 6 dagar eftersom han intehar en etablerad användarbas.
		-- Robert W. Lucky, IEEE President

%
Kom ihåg, UNIX stavat baklänges är Xinu.
		-- Mt.

%
Kom ihåg: använd utloggning logga ut.
		-- Mt.

%
Risch beslut förfarande för integration, inte överraskande,använder en rekursion på antalet och typen av tillägg frånrationella funktioner som behövs för att representera integ. Även omalgoritm följer och kritiskt beror på lämplig strukturav den ingående, såsom i fallet med multivariat faktorisering, kan vi intehävdar att algoritmen är en naturlig. I själva verket, skaparen avdifferential algebra, Ritt, begick självmord i början av 1950-talet,till stor del, hävdas det, eftersom få uppmärksamhet till sitt arbete. Förmodligenhan skulle ha fått mer uppmärksamhet hade han fått algoritmen också.
		-- Joel Moses, "Algorithms and Complexity", ed. J. F. Traub

%
Rad, rad, raden din bitar, försiktigt ner strömmen ...
		-- Joel Moses, "Algorithms and Complexity", ed. J. F. Traub

%
Spara energi: Kör mindre skal.
		-- Joel Moses, "Algorithms and Complexity", ed. J. F. Traub

%
Spara gas, inte använda skalet.
		-- Joel Moses, "Algorithms and Complexity", ed. J. F. Traub

%
Rädda dig själv! Starta i 5 sekunder!
		-- Joel Moses, "Algorithms and Complexity", ed. J. F. Traub

%
Säg "tjugotre-STICK" logga ut.
		-- Joel Moses, "Algorithms and Complexity", ed. J. F. Traub

%
SCCS, källan Motell! Program checka in och aldrig checka ut!
		-- Ken Thompson

%
Vetenskap är att datavetenskap som hydrodynamik är att VVS.
		-- Ken Thompson

%
Forskarna förberedde ett experiment för att ställa den ultimata frågan.De hade arbetat i månader samla en vardera på varje dator som varbyggd. Slutligen den stora dagen var till hands. Alla datorer koppladetillsammans. De ställde frågan, "Finns det en Gud?". lampor börjadeblinkar, blinka och blinkande lite mer. Plötsligt fanns det en högtkrasch, och en blixt kom ned från himlen, slogdatorer, och svetsas alla anslutningar permanent tillsammans. "Detär nu ", kom svaret.
		-- Ken Thompson

%
Scotty: Kapten, vi DIN "kan referera till det!Kirk: Analys, mr Spock?Spock: Kapten, det inte visas i symboltabellen.Kirk: Då är det av yttre ursprung?Spock: Positiv.Kirk: Mr Sulu, går att passera två.Sulu: Aye aye, sir, kommer att passera två.
		-- Ken Thompson

%
"Avsnitt 2.4.3.5 borst (Accept vänta på nya cykel State).I borst AH-funktionen indikerar att den har mottagit enmultimeddelande byte.I borst måste RFD meddelande sändas falska och DAC meddelandemåste skickas passiv sant.AH-funktionen måste avsluta de borst och skriv:(1) ANRS om DAV är falskt(2) AIDS om ATN meddelandet är falskt och varken:(A) grabbarna är aktiv(B) Nor LACS är aktiv "programmerbar Instrumentering
		-- from the IEEE Standard Digital Interface for

%
Säkerhetskontroll: INTRUDER ALERT!
		-- from the IEEE Standard Digital Interface for

%
Verkar dataingenjör, systemvetare och programmerare varpressa ned ett berg när bromsarna gav ut. Skrek de nedberg, allt snabbare, men till slut lyckades sluta att fungera, mer avlycka än något annat, bara inches från tusen droppfot till taggigastenar. Alla fick ut ur bilen:        Den dataingenjör sa, "Jag tror att jag kan fixa det."        System analytiker sade, "Nej, nej, jag tycker att vi borde ta detin till stan och har en specialist titta på det. "        Programmeraren sade, "OK, men först tänker jag att vi ska få tillbakai och se om det gör det igen. "
		-- from the IEEE Standard Digital Interface for

%
SEMINAR MEDDELANDETitel: Är grodor Turing kompatibla?Speaker: Don "The Lion" KnuthSAMMANDRAGFlera forskare vid University of Louisiana har studeratdatorkraft av olika amfibier, grodor i synnerhet. Problemetgroda beräkningsbarhet har blivit en viktig fråga som spänner över alla områdendatavetenskap. Det har visat sig att något beräkningsbar av en amphi-bian gemenskap i en fast storlek damm är beräkningsbar av en groda i samma storlekdamm - det vill säga, grodor är Damm-space komplett. Vi kommer att visa attDet finns en logg-space, polywog-tidsbesparing från någon Turing maskin programtill en groda. Vi kommer att föreslå dessa utgör en riktig delmängd av frog-beräkningsbarfunktioner.Detta är inte bara en låt oss-se-hur-långt-de-grodor-can-jump seminariet.Detta är bara för hardcore amfibie-beräknings människor och deras kollegor.Förfriskningar serveras. Musik spelas.
		-- from the IEEE Standard Digital Interface for

%
Skicka några smutsiga post.
		-- from the IEEE Standard Digital Interface for

%
Sendmail kan vara säkert köra set-användar-id till root.
		-- Eric Allman, "Sendmail Installation Guide"

%
Flera elever ombads att bevisa att alla udda heltal är prime.Den första eleven att försöka göra detta var en mathstudent. "Hmmm ...Brunn, 1 är ett primtal, 3 är ett primtal, 5 är ett primtal, och genom induktion, har vi att allade udda heltal är prime. "Den andra eleven att prova var en man i fysik som kommenterade, "Jag är intesäker på giltigheten av ditt bevis, men jag tror jag ska försöka bevisa det genomexperiment. "Han fortsätter:" Tja, en är utmärkt, 3 är ett primtal, 5 är ett primtal, 7 ärPrime, 9 är ... eh, nio är ... eh, 9 är en experimentell fel, 11 är ett primtal, 13är utmärkt ... Tja, det verkar som du har rätt. "Den tredje elev att prova det var engineering student, som svarade,"Jo, för att vara ärlig, faktiskt, jag är inte säker på svaret heller. Låt ossse ... en är utmärkt, 3 är ett primtal, 5 är ett primtal, 7 är ett primtal, 9 är ... eh, är nio ...Tja, om du närma, är 9 prime, 11 är ett primtal, 13 är ett primtal ... Tja, detverkar rätt. "Inte vara sämre, det datavetenskapliga eleven kommer och säger"Ja, ni två sort've fick rätt idé, men du kommer att hamna tar för lång tid!Jag har bara piskade upp ett program för att verkligen gå och bevisa det. "Han går fram tillsin terminal och kör sitt program. Läsa utgången på skärmen säger han,"1 är ett primtal, en är utmärkt, en är utmärkt, en är utmärkt ..."
		-- Eric Allman, "Sendmail Installation Guide"

%
Hon säljer CSHS av cshore.
		-- Eric Allman, "Sendmail Installation Guide"

%
Shopping på denna grody lilla datorbutik på Galleria för enhelt awwwesome Apple. Fer suuure. Jag menar Äpplen är trevligt du vet?Men, du vet, det är denna söt kille som arbetar där och han säger attVAX s är svalare! Jag menar jag vet inte riktigt, du vet? Han säger att hanhar detta helt tubulär VAX hemma och det är fyllda med minne-to-the-max!Höger, ja. Och han vill ta mig hem för att visa det för mig. Herregud!Jag är suuure. Gag mig med en Prime!
		-- Eric Allman, "Sendmail Installation Guide"

%
Simuleringar är som minikjolar, visar de en hel del och dölja det väsentliga.
		-- Hubert Kirrman

%
skldfjkl jklsR% ^ & (IXDRTYju187pkasdjbasdfbuilh; asvgy8p 23r1vyui 135 2kmxsij90TYDFS $$ b jkzxdjkl bjnk, j nk; <[] [; - == - <<<<< ", [,[Hjioasdvbnuio; buip ^ & (FTSD $% * VYUI: buio; sdf} [asdf ']sdoihjfh (_YU * G & F ^ * CTY98yNu ser vad du har gått och gjort! Du har brutit det!
		-- Hubert Kirrman

%
Långsamt och säkert UNIX kröp upp på Nintendo användare ...
		-- Hubert Kirrman

%
Så du ser Antonio, varför oroa sig för en liten kärna dump, va? I verklighetenalla kärn dumpar händer i samma ögonblick, så kärnan dumpa dig kommer att hai morgon, varför redan hände det. Du ser, det är bara en liten universellrekursiva skämt som trådar våra liv genom den oändliga potentialdet ögonblick. Så somnar, Antonio, kan din tråd bryta helstoch kasta dig ut ur säkra säkerheten i det ögonblick i den mörka tomrumevighet, anti-tiden. Så gå att sova ...
		-- Hubert Kirrman

%
Mjukvara produktionen antas vara en linjefunktion, men det körssom en stabsfunktion.
		-- Paul Licker

%
Mjukvaruleverantörer försöker göra sina programpaket mer"användarvänlig". ... Deras bästa sättet hittills har varit att vidta allagamla broschyrer och stämpla orden "användarvänliga" på omslaget.[Pot. Vattenkokare. Svart.]
		-- Bill Gates, Microsoft, Inc.

%
Några av mina läsare frågar mig vad en "seriell port" är.Svaret är: Jag vet inte.Är det något slags vin du har med frukost?
		-- Bill Gates, Microsoft, Inc.

%
Somliga hävdar att UNIX inlärningskurvan är brant, men åtminstone dubara måste klättra det en gång.
		-- Bill Gates, Microsoft, Inc.

%
Vissa programmeringsspråk lyckas ta till sig förändringar, men tål framsteg.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Någon terminal sjunker bitar. Jag hittade en stapel av dem ihörn.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Något mystiskt bildas, född i den tysta tomrum. Väntarensam och orörlig, är det på en gång stilla och ändå i ständig rörelse. Det ärkällan till alla program. Jag vet inte sitt namn, så jag kommer att kalla detTao of Programming.Om Tao är bra, då operativsystemet är stor. OmOperativsystemet är stor, då kompilatorn är stor. Om kompilatorn ärstörre, då ansökningarna är stor. Användaren är nöjd och det finnsharmoni i världen.Tao av ​​programmering strömmar långt borta och avkastningen på vindmorgon.
		-- Geoffrey James, "The Tao of Programming"

%
På tal som någon som har fördjupat sig i den invecklade PL / I, jag är säker påatt endast Verkliga Män kunde ha skrivit en sådan maskin-hogging, cykel väckande,allomfattande monster. Tilldela en matris och frigöra mellersta tredjedelen?Säker! Varför inte? Multiplicera en teckensträng ibland lite sträng och tilldelaleda till en flottör decimal? Varsågod! Frigöra en reglerad variabel förfarandeparameter och omfördela det innan de passerar den tillbaka? Overlay tre olikatyper av variabel på samma minnesplats? Allt du säger! Skriv enrekursiv makro? Tja, nej, men Real Män använder scanna. Hur kunde ett språkså uppenbart utformade och skriven av verkliga Män inte vara avsedda för Real Man använder?
		-- Geoffrey James, "The Tao of Programming"

%
***** Special AI seminarium (abstract)Det har varit allmänt känt att AI program kräver expertkunskapFör att prestera bra i komplexa domäner. Men enbart kunskap är intetillräckligt för vissa tillämpningar; visdom behövs också. Följaktligen,Vi har utvecklat en ny metod för artificiell intelligens som vi kallar"Visdom engineering". Som ett test av våra idéer, har vi skrivit Immanuel envisdom baserat system för uppgiften domänen i västra filosofiskt tänkande.Immanuel tillfördes initialt med 200 visdomsheter som innehöll visdomom sådana elementära begrepp som sinnet, materia, som, intet, och såvidare. Immanuel tilläts därefter att röra sig fritt, styrs av den heuristiskaregler som ingår i dess heterarchically organiserade meta visdom bas. Immanuellyckats återupptäcka de flesta av de viktiga filosofiska idéer utvecklasi västerländsk kultur under loppet av de senaste 25-talen, inklusive sådanaunderliggande Platons teori regerings Kants metafysik, Nietzsches teorivärde, och Husserls fenomenologi. I detta seminarium kommer vi att beskrivaImmanuel prestationer och intern arkitektur. Vi kommer också kortfattatdiskutera våra senaste ansträngningar att tillämpa visdom teknik till oljeutvinning.
		-- Geoffrey James, "The Tao of Programming"

%
Personalmöte i konferensrummet i% d minuter.
		-- Geoffrey James, "The Tao of Programming"

%
Personalmöte i konferensrummet i 3 minuter.
		-- Geoffrey James, "The Tao of Programming"

%
Standarder är avgörande. Och det bästa med standarder är: det finnsså ____ många att välja mellan!
		-- Geoffrey James, "The Tao of Programming"

%
Fortfarande några buggar i systemet ... Someday jag måste berätta om UncleNahum från Maine, som tillbringade år försöker korsa en manet med en Shadså att han kunde föda benfritt Shad. Sitt experiment misslyckades också, och hanavvecklas med beniga maneter ... som var knappast värt besväret. det finnsmycket liten uppmaning till dem där uppe.
		-- Allucquere R. "Sandy" Stone

%
Snålhet med privilegier är vänlighet i förklädnad.
		-- Guide to VAX/VMS Security, Sep. 1984

%
	Sluta! Den som crosseth bron of Death, måste svara förstdessa frågor tre, innan den andra sidan han se!	"Vad heter du?""Sir Brian Bell.""Vad är ditt uppdrag?""Jag söker den heliga graal.""Vad är fyra gemener som inte är juridiska flagga argumenttill Berkeley UNIX-versionen av `ls '?""Jag, er .... AIIIEEEEEE!"
		-- Guide to VAX/VMS Security, Sep. 1984

%
*** STUDENT FRAMGÅNGAR ***Många av våra elever har gått vidare för att nå stora framgångar inom alla områden avprogrammering. En tidigare student utvecklat begreppet personligbrev. Betyder uttrycket "Dear Mr (ange namn), Du kanske redan vara envinnare !, "låter det bekant? En annan elev skriver" Efter bara fem lektioner jagsålde en "My mest oförglömliga Program" artikeln Frätande Computing magazine.En annan av våra studenter skriver: "Jag har nyligen avslutat en databasadministrationtill min avdelningschef. Mitt program rörde vid honom så djupt att hanvar mållös. Han berättade senare att han aldrig hade sett ett sådant program ihela hans karriär. Tack, berömda Programmerare skola; bara du kundehar gjort detta möjligt. "Skicka för vår inledande broschyr som förklarari vaga detalj driften av den berömda programmerare Skolan, och du kommervara berättigad att vinna en möjlig chans att komma in en ritning, vinnaren somkan tävla om en samling av fria stek knivar. Om du inte gör det nu, kommer du hatarsjälv på morgonen.
		-- Guide to VAX/VMS Security, Sep. 1984

%
Sådana insatser är nästan alltid långsamt, mödosamt, politisk, småaktiga, tråkig,otympligt, otacksam och ytterst kritiskt.
		-- Leonard Kleinrock, on standards efforts

%
Antag för ett ögonblick att bilindustrin hade utvecklats på sammatakt som datorer och under samma period: hur mycket billigare och mereffektivt skulle nuvarande modeller vara? Om du inte redan har hörtAnalogt svaret splittring. Idag skulle du kunna köpa enRolls-Royce för $ 2,75, skulle det göra tre miljoner miles till gallon, ochdet skulle ge tillräckligt med ström för att driva drottning Elizabeth II. Och om duvar intresserade av miniatyrisering, kan du placera ett halvt dussin av dem påett knappnålshuvud.
		-- Christopher Evans

%
Swap läsfel. Du förlorar ditt sinne.
		-- Christopher Evans

%
Syntaktiskt socker orsakar cancer i semikolon.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
System checkpoint komplett.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
System går ner vid 01:45 i eftermiddag för disk kraschar.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
System går ner vid fem i eftermiddag för att installera schemaläggare bugg.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
System går ner i 5 minuter.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
System omstart, vänta ...
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
    *** Avstängning meddelande från rot ***System går ner i 60 sekunder
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Systems har delsystem och delsystem har delsystem och så vidare adoändlighet - det är därför vi alltid börja om från början.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
System programmerare är de höga präster låg kult.
		-- R. S. Barton

%
Testning kan visa pres buggar, men inte deras frånvaro.
		-- Dijkstra

%
Tex är potentiellt den viktigaste uppfinningen i sättning i dettaårhundrade. Det införs ett standardspråk för dator typografi, och itermer av vikt kan rangordna nära införandet av Gutenberg pressen.
		-- Gordon Bell

%
"Textbehandling har gjort det möjligt att höger motivera någon idé, ävenen som inte kan motiveras på någon annan grund. "
		-- J. Finnegan, USC.

%
Det betyder inte beräkna.
		-- J. Finnegan, USC.

%
... Att begreppen "hårdvara", och "programvara" bör förlängas medbegreppet Liveware - är den som producerar programvara för användning påhårdvara. Detta ger en uppenbar utvidgning till begreppet monitorer.En Liveware monitor är en person som ägnar sig åt uppgiften att se till attLiveware inte störa realtidsprocesser, åberoparREALTID bödeln att ta bort Liveware som negativt påverkar ...
		-- Linden and Wihelminalaan

%
"Det är rätt, den versaler skift fungerar bra på skärmen, mende är inte kommer ut på den jävla skrivare ... Håll? Visst, jag ska hålla. "
		-- e.e. cummings last service call

%
Det är det om personer som tror att de hatar datorer. Vad deverkligen hatar är usel programmerare.
		-- Larry Niven and Jerry Pournelle in "Oath of Fealty"

%
"Cutting edge" blir ganska tråkig.
		-- Andy Purshottam

%
11 är för personer med stolthet 10 och plånbok av en åtta.
		-- R. B. Greenberg [referring to PDPs?]

%
Frånvaron av etiketter [i ECL] är förmodligen en bra sak.
		-- T. Cheatham

%
Algoritmen för att finna den längsta bana i en graf är NP-fullständigt.För dig system människor, innebär att det är * väldigt långsamt *.
		-- Bart Miller

%
"Algoritmen att göra det är extremt otrevlig. Du kanske vill rånanågon med det. "
		-- M. Devine, Computer Science 340

%
Analytical Engine väver algebraiska mönster precis som Jacquardvävstol väver blommor och blad.
		-- Ada Augusta, Countess of Lovelace, the first programmer

%
"Den dåliga rykte UNIX har fått är helt oförtjänt, som på av människorsom inte förstår, som inte har kommit in där och försökte något. "
		-- Jim Joyce, owner of Jim Joyce's UNIX Bookstore

%
Öl kylda dator inte skadar ozonskiktet.[Om jag kan läsa mina anteckningar från Be Dr. Mike session på Baycon, jagtror han tillade att ölet kylda dator använder "Forget EndastMinne ". Ed.]
		-- John M. Ford, a.k.a. Dr. Mike

%
Den bästa boken om programmering för en lekman är "Alice i Underlandet";men det beror på att det är den bästa bok om något för en lekman.
		-- John M. Ford, a.k.a. Dr. Mike

%
Det bästa sättet att påskynda en Macintoy är 9,8 meter per sekund per sekund.
		-- John M. Ford, a.k.a. Dr. Mike

%
Den bogosity meter bara knuten.
		-- John M. Ford, a.k.a. Dr. Mike

%
Buddha, Gudomen, bosatt riktigt lika bekvämt i kretsarna i endigital dator eller redskap med en cykel överföring som han gör på toppenav ett berg eller i kronbladen på en blomma. Att tro något annat är att förnedraBuddha - vilket är att förnedra sig själv.
		-- Robert Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
De fel som du måste undvika är de som ger användaren inte barabenägenheten att få på ett plan, men också tiden.
		-- Kay Bostic

%
"The C Programming Language - Ett språk som kombinerar flexibiliteten hosassembler med kraften av assembler. "
		-- Kay Bostic

%
Kläderna har ingen kejsare.
		-- C. A. R. Hoare, commenting on ADA.

%
Datorindustrin är journalister i 20-årsåldern som står i vördnad förföretagare i sina 30-talet som anställer säljare i deras 40-talet och50 och betala dem i 60- och 70-talet för att få sin marknadsföring i80-talet.
		-- Marty Winston

%
Datorn är att informationsindustrin ungefär vadcentral kraftstation är att den elektriska industrin.
		-- Peter Drucker

%
"Computer fick mig att göra det."
		-- Peter Drucker

%
Beräknings fältet är alltid i behov av nya klichéer.
		-- Alan Perlis

%
Sambandet mellan det språk som tror att vi / program och de problemoch lösningar som vi kan föreställa oss är mycket nära. Av denna anledning begränsandespråkfunktioner med avsikten att eliminera programmerare fel är i bästa fallfarlig.
		-- Bjarne Stroustrup

%
Dag till dag travails av IBM programmerare är så roligt att de flesta avoss som har turen att aldrig ha varit en - som att seCharlie Chaplin försöker laga en sko.
		-- Bjarne Stroustrup

%
Debatten rasar på: Är PL / I Bachtrian eller dromedar?
		-- Bjarne Stroustrup

%
Skillnaden mellan konst och vetenskap är att vetenskapen är vad viförstår tillräckligt bra för att förklara för en dator. Konst är allt annat.
		-- Donald Knuth, "Discover"

%
Skivorna blir fullt; rensa en fil idag.
		-- Donald Knuth, "Discover"

%
"Den elfte budet var` Du skall Compute 'eller' Du skall ickeBeräkna "- jag glömmer vilken".
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Sätta in vägleder till nordamerikanska HANARARTER: Cranial MänUnderarter: The Hacker (homo computatis)Uppvaktning & Mating:På grund av extrem fattigdom, HOMO COMPUTATIS upprätthåller en nära evigtillstånd av sexuell beredskap. Parningsbeteende alternerar mellanbesvärliga blyghet och plötsliga framsteg. När han till slut kompisar, hanväljer en kvinnlig ingenjör med en unblinking stare, en stram mun, ochen komplett samling av Campbells soppa-burk recept.Spåra:Soptunnor full av ljusgrönt och vitt perforerat papper och gamlakopior av Allen-Bradley katalog.kommentarer:Extremt förtjust i dåliga vitsar och skämt som behöver långa förklaringar.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Sätta in vägleder till nordamerikanska HANARARTER: Cranial MänUnderarter: The Hacker (homo computatis)Beskrivning:Gängliga och svaga, har hackaren en hög panna och gallring hår.Chef oproportionerligt stor och krokig framåt, hy glåmig ochsightly grå från CRT belysning. Han har tunga svarta glasögonoch en blick av intensiv koncentration, vilken kan bero på en programvaraproblem eller till en fläsk-och-bönor frukost.ludd:HOMO COMPUTATIS såg en Brylcreem annons femton år sedan och trodde det.Följaktligen är crest smord ner, med undantag för den cowlick.Låt:En ganska klagande "Är det?"
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Sätta in vägleder till nordamerikanska HANARARTER: Cranial MänUnderarter: The Hacker (homo computatis)fjäderdräkt:Alla kläder har en något skrynklig ser ut som om de kom fråntoppen av tvättkorgen. Style varierar med status. hacker cheferbära grå polyester byxor, rosa eller pastell skjortor med breda kragar,och paisley band; Personalen bär fastsatt upp baggy manchester byxor, viteller blå skjortor med button-down kragar och pennhållare i fickan.Både chefer och personalen bära löparskor att arbeta, och en svartplast digital klocka med miniräknare.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Första gången är det en kludge!Den andra, ett trick.Senare, det är en väl etablerad teknik!
		-- Mike Broido, Intermetrics

%
Den första versionen alltid får kastas bort.
		-- Mike Broido, Intermetrics

%
Flödesschemat är en mest grundligt översåld bit av programdokumentationen.
		-- Frederick Brooks, "The Mythical Man Month"

%
Följande citat är från sidan 4-27 av MSCP enkel disk funktionerHandbok som är en del av manualer UDA50 Programmerare Doc Kit:Såsom angivits ovan, är värd cirkelns area strukturerad som en vektor avlogiska block. Ur prestandasynpunkt, är det emellertid merlämpligt att visa värdområdet som fyrdimensionell hyper-kuben,fyra dimensioner är cylinder, grupp, spår och sektor.. . .Med hänvisning till vår hyper-kub analogi, uppsättningen av potentiellt tillgängligablock bildar en linje parallell med körbanans axel. Denna linje flyttarparallellt med sektoraxeln, linda runt när den når kantenav hyperkuben.
		-- Frederick Brooks, "The Mythical Man Month"

%
Fontänen koden har skärpts något så att du inte längre kan doppaobjekt i en fontän eller dricka från en medan du svävar i luftenpå grund av levitation.Teleportera till helvetet via en teleporte fälla kommer inte längre att skeom tecknet inte har brandmotstånd.
		-- README file from the NetHack game

%
Målet för datavetenskap är att bygga något som kommer att pågå istone tills vi har byggt färdigt den.
		-- README file from the NetHack game

%
Gurus Unix Meeting of Minds (Gumm) sker onsdag april1, 2076 (se det i din evighetskalender program), 14 fot ovanmarken direkt framför Milpitas Gumps. Medlemmarna kommer grepvarandra vid handen (efter intro), yacc mycket, rök filtreradeschroots i rör, chown med gafflar, använda wc (såvida uuclean), fseektrevliga zombie processer, band, och sova, men inte, hoppas vi, OD. Tredagar kommer att ägnas åt diskussion om konsekvenserna av whodo. Tvåsekunder har tilldelats för en fullständig genomgång av alla användarvänliga funktioner av Unix. Seminarier inkluderar "allt du vet ärFel ", som leds av Tom Kempson," Batman eller katt: man "leds av Richie Dennis?"Cc C? Si! Si!" ledd av Kerwin Bernighan och "Dokument Unix, är duSkojar? "Under ledning av Jan Yeats. Ingen Reader service No. är nödvändigt eftersomalla GUGUs (Gurus Unix grupp användare) redan vet allt vikunde berätta.
		-- "Get GUMMed," Dr. Dobb's Journal, June '84

%
Killen på höger Inte en chansKillen till höger har Osborne 1, en fullt fungerande datorsystemi ett bärbart paket storleken på en portfölj. Killen till vänster har enUzi kulsprutepistol dold i sin attachéväska. Även i fallet är fyrafullastad, 32-runda klipp med 125-korn 9mm ammunition. Ägaren avUzi kommer att få mer taktiska eldkraft levereras - och levereras irikta - på kortare tid, och med mindre ansträngning. Allt för $ 795. Det är oundvikligt.Om du går upp mot en kille med en Osborne 1 - eller någon personligdator - han är den som har problem. En runda från en Uzi kan zipgenom tio inches av massiv furu trä, så kan ni föreställa er vad det kommer att göratill strukturskum akryl och aluminiumplåt. I själva verket, löstagbara tidningarför Uzi finns i 25-, 32-, och 40-runda kapacitet så att du kanta ut ett helt kontor full av Apple II eller IBM Personal Computers bundnai Ethernet eller andra nätverk lokala området. Vad om den nya 16-bitarsdatorer, som Lisa och Fortune? Även med Winchester backup,De är ingen match för Uzi. En snabb burst och de kommer att ta reda på vadUnix betyder. Gör din befäl stolt. Få en Uzi - och komma hemen vinnare i kampen för kontorsautomatvapen.
		-- "InfoWorld", June, 1984

%
Den mänskliga hjärnan fungerar normalt endast tio procent av sin kapacitet- Resten är overhead för operativsystemet.
		-- Nicholas Ambrose

%
IBM 2250 är imponerande ...om man jämför med ett system försäljning för en tiondel sitt pris.
		-- D. Cohen

%
IBM förvärv av ROLM ger ny innebörd åt uttrycket "twisted pair".
		-- Howard Anderson, "Yankee Group"

%
Tanken att en godtycklig naiv människa ska kunna korrekt använda en vissverktyg utan utbildning eller förståelse är ännu mer fel för beräkning ändet är för andra verktyg (t ex bilar, flygplan, vapen, motorsågar).
		-- Doug Gwyn

%
Den sista gången någon sa, "Jag tycker jag kan skriva mycket bättre med ett ordprocessor. ", svarade jag," De brukade säga samma sak om droger. "
		-- Roy Blount, Jr.

%
Ju mindre tid planering, desto mer tid programmering.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 10: ENKELSIMPLE är en akronym för Sheer Idiot Monopurpose programmeringsspråkMiljö. Detta språk, som utvecklats vid Hannover College förTekniska Misfits, har utformats för att göra det omöjligt att skriva kodmed fel i det. Uttalandena är därför begränsad till Begin,END och STOP. Oavsett hur du ordnar uttalanden, kan du inte göraett syntaxfel. Program skrivna i SIMPLE göra något användbart. Såledesde uppnå de resultat av program skrivna i andra språk utandet tråkiga, frustrerande processen för testning och felsökning.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 12: LITHPDetta annars utmärker språk kännetecknas av avsaknad avett "S" i sin teckenuppsättning; användare måste ersätta "TH". LITHP sägsvara användbara vid protheththing lithtth.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 13: SlobolSlobol är mest känd för hastighet, eller avsaknaden av den, av dess kompilator.Även om många kompilatorer kan du ta en fika medan desammanställa, Slobol kompilatorer kan du resa till Bolivia för att plockakaffe. Fyrtiotre programmerare är kända för att ha dött av tristesssitter vid sina terminaler i väntan på en Slobol programsammanställa. Trötta Slobol programmerare vänder sig ofta till en närstående (menoändligt snabbare) språk, kokain.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 14 - VALGOLVALGOL njuter en dramatisk ökning av popularitet överindustri. VALGOL kommandon inkluderar verkligen, som, ja, och Y * veta.Variabler tilldelas med = LIKE och = Helt operatörer. Andraoperatörer inkluderar "California booleska", AX och NOWAY. slingor äruppnås med FOR SURE konstruera. Ett enkelt exempel:LIKE, Y * VETA (jag menar) STARTIF PIZZA = LIKE Bitchen OCHGUY = LIKE rörelement ochDalflickan = LIKE Grody ** MAX (FERSURE) ** 2DÅFör i = LIKNANDE en TILL OH * KANSKE 100DO * WAH - (DIKT ** 2); BARF (I) = helt brutto (OUT)		SÄKERLIKE, BAG detta program, VERKLIGEN; LIKE TOTALT (Y * vet); JAG ÄR SÄKER	GÅ TILL KÖPCENTRETVALGOL kännetecknas också av sin ovänliga felmeddelanden. Förexempel, när användaren gör ett syntaxfel visar tolkenmeddelande Gag mig med en sked! En framgångsrik compile kan benämnas maximaltGRYMT BRA!
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 15 - DogoUtvecklat vid Massachusetts Institute of lydnadsträning, DOGODOGO inleder en ny era av datorkunnig husdjur. Dogo kommandon inkluderarSIT, stanna, fot, och rulla över. Ett innovativt inslag i DOGO är "valpgrafik ", en liten cocker spaniel som ibland lämnar en deposition somden färdas över skärmen.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 16: C-Detta språk namngavs för betyget emot av dess skapare, då hanlade fram det som ett klassprojekt i en examen programmerings klass. C- är bästbeskrivs som ett programmeringsspråk "låg nivå". I själva verket, det språki allmänhet kräver mer C- uttalanden än maskin kod uttalandenutföra en given uppgift. I detta avseende är det mycket lik COBOL.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 17: SARTREUppkallad efter den sena existentiella filosofen, är SARTRE en extremtostrukturerad språk. Uttalanden i SARTRE har något syfte; de bara är.Således SARTRE program kvar att definiera sina egna funktioner. SARTREprogrammerare tenderar att vara tråkig och deprimerad, och är inget kul på fester.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 18: FemteFEMTE är en precisions matematiskt språk som datatypernahänvisa till kvantiteten. Datatyperna varierar från CC, uns, SHOT, ochMANICK till femte (därav namnet på det språk) liter, MAGNUM ochBLOTTO. Kommandon hänvisar till ingredienser såsom Chablis, Chardonnay,CABERNET, gin, vermouth VODKA, SCOTCH och WHATEVERSAROUND.De många versioner av den femte språket speglar den sofistikerade ochfinansiella ställning av dess användare. Kommandon i ELITE dialekt inkluderarVSOP och LAFITE, medan kommandon i rännstenen dialekt inkluderar Hootchoch rippel. Det senare är en favorit av frustrerade FRAMÅT programmeraresom sluta använda detta språk.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 2: RenéUppkallad efter den berömda franska filosofen och matematikern René Descartes,RENE är ett språk som används för artificiell intelligens. Språket ärutvecklats vid Chicago Center of Machine Politik och programmering under enbevilja från Jane Byrne Victory Fund. En talesman beskrev språksom "lika stor som dis [sic] staden vår."Centret är mycket nöjd med utvecklingen hittills. De säger att de har nästanlyckats få en VAX att tänka. Men källor inne iorganisation säga att varje gång maskinen inte tror att det upphör att existera.
		-- Roy Blount, Jr.

%
De mindre kända programmeringsspråk # 8: LaidbackDetta språk utvecklades i Marin County Center för T'ai Chi,Vekhet och Programmerings (nu nedlagda), som ett alternativ tillmer intensiv atmosfär i närheten Silicon Valley.Centret var perfekt för programmerare som velat dra i badtunnor medande arbetade. Tyvärr få programmerare kunde överleva där eftersomcentrum förbjöd Pizza och Coca-Cola till förmån för Tofu och Perrier.Många sörjer nedläggningen av Laidback på grund av sitt rykte som en mild ochicke-hotande språk eftersom alla felmeddelanden är i gemener. FörExempelvis svarade Laidback till syntaxfel med budskapet:"Jag hatar att störa dig, men jag bara inte kan relatera till det. Kandu hitta tid att prova igen? "
		-- Roy Blount, Jr.

%
Macintosh är Xerox teknik som bäst.
		-- Roy Blount, Jr.

%
Trollkarlen Elfenbenstornet tog sin senaste uppfinning förMaster programmerare att undersöka. Magikern hjul en stor svart låda imästare kontor medan befälhavaren väntade under tystnad."Detta är en integrerad, distribueras, allmänt ändamål arbetsstation"började trollkarlen "ergonomiskt utformad med en egen driftssystemet, sjätte generationens språk, och flera toppmoderna användargränssnitt. Det tog mina assistenter flera hundra manår att bygga.Är det inte fantastiskt? "Befälhavaren höjde ögonbrynen en aning. "Det är verkligen häpnadsväckande," hansa."Corporate högkvarter har befallt", fortsatte trollkarlen "somalla använder denna arbetsstation som en plattform för nya program. Håller du medtill detta?""Visst", svarade befälhavaren, "Jag kommer att få det transporteras tilldatacenter omedelbart! "Och trollkarlen återvände till sitt torn, välnöjd.Flera dagar senare, vandrade en novis i kontoret av befälhavarenprogrammerare och sa, "Jag kan inte hitta notering för mitt nya program. Hardu vet var det kan vara? ""Ja", svarade befälhavaren "listor staplas på plattformeni datacentret. "
		-- Geoffrey James, "The Tao of Programming"

%
Master programmerare flyttar från program till program utan rädsla. Nejförändring i förvaltningen kan skada honom. Han kommer inte att avfyras, även om projektetavbryts. Varför är detta? Han är fylld med Tao.
		-- Geoffrey James, "The Tao of Programming"

%
Köttet är ruttet, men spriten håller ut.Computer översättning av "Anden är villig, men köttet är svagt."
		-- Geoffrey James, "The Tao of Programming"

%
Meta-Turingtestet räknas en sak som intelligent om det syftar till attutforma och tillämpa turingtest till föremål för sin egen skapelse.
		-- Lew Mammel, Jr.

%
Den misnaming av ämnesområden är så vanligt som leder till vad som kan varaallmänna system lagar. Till exempel, Frank Harary föreslog en gång den lag somnågot fält som hade ordet "vetenskap" i sitt namn garanterades därigenominte att vara en vetenskap. Han skulle nämner som exempel militärbranschen, bibliotekScience, statsvetenskap, Hemkunskap vetenskap, samhällsvetenskap, och datorVetenskap. Diskutera allmän av denna lag, och möjliga orsaker till dessprognosförmåga.tänkande "
		-- Gerald Weinberg, "An Introduction to General Systems

%
Ju mer data jag stämpla i detta kort, desto ljusare blir, ochsänka utskick kostnad.
		-- S. Kelly-Bootle, "The Devil's DP Dictionary"

%
Den viktigaste tidig produkt på väg att utveckla en bra produktär en ofullkomlig version.
		-- S. Kelly-Bootle, "The Devil's DP Dictionary"

%
Den rörliga markören skriver, och efter att ha skrivit, blinkar.
		-- S. Kelly-Bootle, "The Devil's DP Dictionary"

%
Nätet är som ett stort hav av lutfisk med små dinosaurier hjärnor inbäddadei det här och där. Varje given sked kommer troligen att ha en IQ på en, menenstaka skedar kan ha en IQ mer än sex gånger så!
		-- James 'Kibo' Parry

%
Nya testamentet ger grunden för modern dator kodningsteori,i form av en bekräftelse av det binära talsystemet.Men låt din kommunikation vara ja, ja; nej, nej:för allt som är mer än av ondo.
		-- Matthew 5:37

%
Nästa person att nämna spaghetti staplar för mig kommer att hahuvudet knackade bort.
		-- Bill Conrad

%
Det fina med standarder är att det finns så många av dem att välja mellan.
		-- Andrew S. Tanenbaum

%
Det trevligaste Alto är att det inte köra snabbare på natten.
		-- Andrew S. Tanenbaum

%
Föreställningen om en "record" är en föråldrad kvarleva av dagarna i 80-kolonnkort.
		-- Dennis M. Ritchie

%
Antalet argument är oviktigt om inte en del av dem är korrekta.
		-- Ralph Hartley

%
Antalet datavetare i ett rum är omvänt proportionelltill det antal fel i sin kod.
		-- Ralph Hartley

%
Antalet UNIX installationer har vuxit till 10, med mer väntat.
		-- The Unix Programmer's Manual, 2nd Edition, June 1972

%
Den enda skillnaden mellan en bilförsäljare och en dator försäljare äratt bilförsäljare vet att han ljuger.
		-- The Unix Programmer's Manual, 2nd Edition, June 1972

%
Det enda billigare än hårdvara talas.
		-- The Unix Programmer's Manual, 2nd Edition, June 1972

%
Det enda som är värre än X Windows: (X Windows) - X
		-- The Unix Programmer's Manual, 2nd Edition, June 1972

%
Partiet skjuts upp till en bubbelpool, ja. Fullt påklädd, kan jag tillägga.
		-- IBM employee, testifying in California State Supreme Court

%
Den personliga datorn marknaden är ungefär lika stor som den totala potatischipsmarknadsföra. Nästa år kommer det att vara ungefär hälften så stor som sällskapsdjur livsmedelsmarknaden ochnärmar sig snabbt den totala försäljningen av strumpbyxor världen "
		-- James Finke, Commodore Int'l Ltd., 1982

%
Den primära funktionen för konstruktören är att göra sakersvårt för tillverkaren och omöjligt för servicemannen.
		-- James Finke, Commodore Int'l Ltd., 1982

%
Det primära syftet med DATA uttalande är att ge namn åt konstanter;i stället för att hänvisa till pi som 3,141592653589793 vid varje utseende,variabel PI kan ges detta värde med en DATA uttalande och används i ställetav den längre formen av det konstanta. Detta förenklar också modifieraprogram, bör värdet av pi förändring.
		-- FORTRAN manual for Xerox Computers

%
Problemet med ingenjörer är att de tenderar att fuska för attfå resultat.Problemet med matematiker är att de tenderar att arbeta på leksakenproblem för att få resultat.Problemet med program kontrollörer är att de tenderar att fuska vidleksak problem för att få resultat.
		-- FORTRAN manual for Xerox Computers

%
Problemen företagsekonomi i allmänhet och databashantering isynnerhet är mycket svårt för människor som tror på IBMese, sammansattamed slarviga engelska.
		-- Edsger Dijkstra

%
Programmet är inte debuggade till sista användaren är död.
		-- Edsger Dijkstra

%
Programmerarna gamla var mystisk och djup. Vi kan inte förståderas tankar, så allt vi gör är att beskriva deras utseende.Aware, som en räv passerar vattnet. Alert, som en allmän påslagfält. Kind, som en värdinna hälsning sina gäster. Enkelt, som uncarvedblock av trä. Ogenomskinlig, som svarta pooler i mörka grottor.Vem kan berätta hemligheter deras hjärtan och sinnen?Svaret finns endast i Tao.
		-- Geoffrey James, "The Tao of Programming"

%
Beviset att IBM uppfann inte bilen är att den har en rattoch en accelerator i stället för sporrar och rep, för att vara förenliga med en häst.
		-- Jac Goudsmit

%
Anledningen datachips är så små är datorer inte äter mycket.
		-- Jac Goudsmit

%
Den relativa betydelsen av filer beror på deras kostnad i form av denmänsklig ansträngning som krävs för att regenerera dem.
		-- T. A. Dolotta

%
Vägen till helvetet är stenlagd med NAND-grindar.
		-- J. Gooding

%
Försäljaren och systemanalytiker tog fart för att tillbringa en helg iskog, jakt björn. De hade hyrt en stuga, och när de kom dit, togsina ryggsäckar och sätta dem inne. Vid vilken punkt vände säljaretill sin vän, och sa, "du packar medan jag gå och hitta oss en björn."Förbryllad, avslutade analytikern uppackning och sedan gick och satte sigpå verandan. Snart kunde han höra prasslande ljud i skogen. ljudenfick närmare - och högre - och plötsligt fanns försäljare, kör somhelvete över clearing mot kabinen, förföljd av en av de största ochmest våldsamma grizzly bär analytikern hade någonsin sett."Öppna dörren!", Skrek försäljaren.Analytikern vispad öppna dörren, och försäljaren sprang till dörren,plötsligt stannade och steg åt sidan. Björnen, oförmögen att stoppa, fortsattegenom dörren och in i kabinen. Försäljaren smällde igen dörren stängdoch flinade på sin vän. "Fick honom!", Utropade han, "nu, din hud dettaen och jag ska gå prassla oss upp en annan! "
		-- J. Gooding

%
Sendmail Konfigurationsfilen är en av de filer som ser ut som någonslå huvudet på tangentbordet. Efter att ha arbetat med det ... jag kan se varför!
		-- Harry Skelton

%
Den så kallade "stationära metafor" av dagens arbetsstationer är istället en"Flygplan-sits" metafor. Den som har blandas en mantel full av pappernär du sitter mellan två portly passagerare kommer att känna igen skillnaden -kan man se endast en mycket få saker på en gång.
		-- Fred Brooks

%
Steady state diskar är full.
		-- Ken Thompson

%
Systemet var nere för säkerhetskopior från 05:00 till 10:00 i lördags.
		-- Ken Thompson

%
Systemet kommer att vara nere i 10 dagar för förebyggande underhåll.
		-- Ken Thompson

%
Tao tar inte sidor;Det ger upphov till både vinster och förluster.Guru inte ta ställning;Hon välkomnar både hackare och lusers.Tao är som en stack:data ändras men inte strukturen.ju mer du använder den, desto djupare blir;ju mer man talar om det, desto mindre förstår.Håll i roten.
		-- Ken Thompson

%
Tao är som en glob mönster:begagnad men aldrig använt upp.Det är som extern tomrum:fylld med oändliga möjligheter.Det är maskerat men alltid närvarande.Jag vet inte vem som byggde det.Det kom innan den första kärnan.
		-- Ken Thompson

%
Tao som kan vara tjära (1) edär inte hela Tao.Den väg som kan angesär inte den fullständiga sökvägen.Vi förklarar namnenav alla variabler och funktioner.Ändå Tao har ingen typ specificerare.Dynamiskt bindande, inser du det magiska.Statiskt bindande, du ser bara hierarkin.Ändå magi och hierarkihärrör från samma källa,och denna källa har en nollpekare.Hänvisnings NULL inom NULL,Det är inkörsporten till all trolldom.
		-- Ken Thompson

%
Problemet med datorer är att de gör vad du tala om för dem, inte vaddu vill.
		-- D. Cohen

%
UNIX filosofi innebär i princip ger dig tillräckligt repethänga själv. Och sedan ett par fötter, bara för att vara säker.
		-- D. Cohen

%
Användningen av antropomorf terminologi när man behandlar datorsystemär ett symptom på professionell omognad.
		-- Edsger Dijkstra

%
Användningen av COBOL lamslår sinnet; sin undervisning bör därför varabetraktas som ett brott.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
Värdet av ett program är proportionell mot vikten av sin produktion.
		-- Edsger W. Dijkstra, SIGPLAN Notices, Volume 17, Number 5

%
Den vise programmerare berättas om Tao och följer det. Genomsnittetprogrammerare berättas om Tao och söker efter den. Dåren programmerareberättas om Tao och skrattar åt det. Om det inte vore för skratt, detskulle finnas någon Tao.De högsta ljud är svårast att höra. Framöver är ett sätt attreträtt. Större talang visar sig sent i livet. Även en perfekt programfortfarande har buggar.
		-- Geoffrey James, "The Tao of Programming"

%
Arbetet [mjukvaruutveckling] blir mycket lättare (dvs verktygenvi använder arbete på en högre nivå, mer bort från maskinen, periferoch operativsystem imperativ) än den var för tjugo år sedan, och eftersomav detta, kan kännedom om de interna delarna av ett system blir mindre tillgängliga.Vi kanske kan gräva djupare hål, men om vi inte vet hur man bygger högrestegar, hade vi bästa hopp om att det inte regnar mycket.
		-- Paul Licker

%
Världen går mot sitt slut ... Spara BUFFERTAR !!!
		-- Paul Licker

%
Världen går mot sitt slut. Vänligen logga ut.
		-- Paul Licker

%
Världen är inte oktala trots december
		-- Paul Licker

%
Världen kommer att avslutas under 5 minuter. Logga ut.
		-- Paul Licker

%
Den unga damen hade en ovanlig lista,Kopplat delvis en strukturell svaghet.Hon sätter inga förutsättningar.
		-- Paul Licker

%
THEGODDESSOFTHENETHASTWISTINGFINGERSANDHERVOICEISLIKEAJAVELININTHENIGHTDUDE
		-- Paul Licker

%
... Finns det omkring 5000 personer som ingår i denna kommitté. dessa killarhar svårt att reda ut vad dag för att träffa, och om att äta croissantereller munkar till frukost - att inte tala om hur man definierar hur alla dessa komplexaskikt som kommer att komma överens om.
		-- Craig Burton of Novell, Network World

%
Det finns aldrig några fel som du inte har hittat ännu.
		-- Craig Burton of Novell, Network World

%
Det finns nya meddelanden.
		-- Craig Burton of Novell, Network World

%
Det finns inga spel på detta system.
		-- Craig Burton of Novell, Network World

%
Det kör jobb. Varför går du inte jaga dem?
		-- Craig Burton of Novell, Network World

%
Det finns tre typer av människor: män, kvinnor, och Unix.
		-- Craig Burton of Novell, Network World

%
Det finns tre möjligheter: Pioneers solpanel har vänt sig bort frånsolen; Det finns en stor meteor blockerar transmission; någon laddad StarTrek 3,2 i vår videoprocessor.
		-- Craig Burton of Novell, Network World

%
Det finns två stora produkter som kommer ut ur Berkeley: LSD och UNIX.Vi tror inte att det är en tillfällighet.
		-- Jeremy S. Anderson

%
Det finns två sätt att konstruera en programvara design. Ett sätt är att göradet så enkelt att det inte är självfallet inga brister och den andra är attgöra det så komplicerat att det inte finns några uppenbara brister.
		-- C. A. R. Hoare

%
Det finns två sätt att skriva program felfria; endast den tredje fungerar.
		-- C. A. R. Hoare

%
Det har också varit en del arbete för att tillåta intressant användning av makronamn.Till exempel, om du ville alla dina "creat ()" samtal för att inkludera läsabehörigheter för alla, kan man säga#define creat (fil, mode) creat (fil, mode | 0444)Jag rekommenderar mot denna typ av sak i allmänhet, eftersom detdöljer de förändrade semantiken för "creat ()" i ett makro, potentiellt långt bortafrån dess användningsområden.För att tillåta denna användning av makron, använder förprocessorn en process somär värt att beskriva, om av någon annan anledning än att vi får använda en avde mera roande termer introduceras i C lexikon. Medan ett makro ärbyggs ut, är det tillfälligt odefinierad och en upprepning av makrotNamnet "målad blå" - jag ungen du inte, är detta den officiella terminologi- Så att i framtida genomsökningar av texten makrot kommer inte att utökasrekursivt. (Jag vet inte varför den blå färgen valdes, jag är säker på att detvar resultatet av en lång debatt, spridda över flera möten.)
		-- From Ken Arnold's "C Advisor" column in Unix Review

%
Det finns ingen anledning för varje person att ha en dator i sitt hem.Konvention World Future Society, i Boston, 1977
		-- Ken Olsen (President of Digital Equipment Corporation),

%
Det finns ingen skillnad mellan någon AI program och vissa existerande spel.
		-- Ken Olsen (President of Digital Equipment Corporation),

%
Det var en gång en man som gick till en dator mässa. Varje dag somhan kom in, mannen berättade vakten vid dörren:"Jag är en stor tjuv, känd för mina bedrifter av snatteri. Varvarnat för denna mässa får inte undkomma unplundered. "Detta tal störd vakten kraftigt, eftersom det fanns miljonerdollar av datorutrustning inne, så han såg mannen noggrant.Men mannen bara vandrade från monter till monter, nynnar tyst för sig själv.När mannen lämnade tog vakten honom åt sidan och sökte sina kläder,men ingenting stod att finna.Nästa dag på mässan, återvände mannen och bannade denvakta säger: "Jag flydde med en stor byte igår, men idag kommer att bli ännubättre. "Så vakten såg honom allt tätare, men till ingen nytta.Den sista dagen av mässan, kan vakten hålla sinnyfikenhet inte längre. "Sir Thief", sade han, "jag är så förbryllad, kan jag inte levai fred. Vänligen upplysa mig. Vad är det som du stjäl? "Mannen log. "Jag stjäla idéer", sade han.
		-- Geoffrey James, "The Tao of Programming"

%
Det var en gång en mästare programmerare som skrev ostrukturerade program.En nybörjare programmerare, försöker imitera honom, började också att skriva ostruktureradprogram. När nybörjare bad befälhavaren att utvärdera hans framsteg,herre kritiserade honom för att skriva ostrukturerade program, säger: "Vad ärlämplig för befälhavaren inte är lämplig för nybörjare. Du måsteförstå Tao innan vinna struktur. "
		-- Geoffrey James, "The Tao of Programming"

%
Det var en gång en programmerare som var knuten till domstolen i denwarlord av Wu. Krigsherren frågade programmeraren: "Vilket är lättare att utforma:en redovisning paket eller ett operativsystem? ""Ett operativsystem", svarade programmeraren.Krigsherren yttrade ett utrop av misstro. "Säkert enredovisning paket är trivialt bredvid komplexiteten av ett operativsystemsystemet ", sade han."Inte så", sade programmeraren "när man utformar en redovisning paket,programmeraren fungerar som en medlare mellan människor med olika idéer:hur det ska fungera, hur dess rapporter ska visas och hur det måste överensstämma medskattelagstiftningen. Däremot är ett operativsystem inte begränsat min utanförutseenden. Vid utformningen av ett operativsystem, programmeraren sökerenklaste harmoni mellan maskinen och idéer. Detta är anledningen till att ett operativsystemär lättare att utforma. "Krigsherren Wu nickade och log. "Det är allt bra och väl, mensom är lättare att felsöka? "Programmeraren gjorde inget svar.
		-- Geoffrey James, "The Tao of Programming"

%
Det var en gång en programmerare som arbetade på mikroprocessorer. "Titta påhur bra jag är här ", sade han till en stordator programmerare som kom på besök,"Jag har mitt eget operativsystem och fil lagringsenhet. Jag behöver intedela mina resurser med någon. Programvaran är fristående ochlätt att använda. Varför inte sluta ditt nuvarande jobb och gå med mig här? "Stordator programmerare började sedan att beskriva sitt system till sinvän, säger: "Den stordator sitter som en gammal salvia mediterar imitt i datacentret. Dess hårddiskar ligger end-to-end som en stor oceanav maskiner. Programvaran är en mångfacetterad som en diamant och så inveckladsom en urtida djungel. Programmen, varje unik, rör sig genom systemetsom en snabb-strömmande flod. Det är därför jag är glad där jag är. "Mikrodatorn programmerare, när han hörde detta, tystnade. Mentvå programmerare förblev vänner till slutet av sina dagar.
		-- Geoffrey James, "The Tao of Programming"

%
Det fanns, det dök upp, en mystisk rit om inledande genom vilken,på ett eller annat sätt, nästan varje medlem i teamet passerat. Termenatt de gamla händer som används för denna rit - West uppfann sikt intepraxis - var `registrerar dig". Genom att registrera dig för projektet som du kommit överensatt göra vad som var nödvändigt för att lyckas. Du gick med på att överge, omnödvändiga, familj, fritidsintressen och vänner - om du hade någon av dessa kvar(Och du kanske inte, om du hade skrivit för många gånger tidigare).
		-- Tracy Kidder, "The Soul of a New Machine"

%
Det måste vara mer i livet än sammanställa-and-go.
		-- Tracy Kidder, "The Soul of a New Machine"

%
De kallas datorer helt enkelt eftersom beräkningen är den enda betydandejobb som hittills getts till dem.
		-- Tracy Kidder, "The Soul of a New Machine"

%
De är relativt bra men helt fruktansvärt.
		-- Alan Kay, commenting on Apollos

%
De verkar ha lärt sig vanan att huka inför auktoritet även närfaktiskt inte hotad. Hur mycket trevligt för myndigheten. Jag beslutade att intelära denna läxa.
		-- Richard Stallman

%
Tänk på det! Med VLSI kan vi packa 100 ENIACs i 1 kvm. Cm.!
		-- Richard Stallman

%
Tänk på din familj i kväll. Försök att krypa hem efter att datorn kraschar.
		-- Richard Stallman

%
Denna "brain-skadade" epitetet blir i högsta grad överarbetad. När vi kantala om någon eller något är bristfällig, nedsatt, fördärvad, bortskämd;batty, GALEN, bonkers, buggy, knäckt, galen, gök, tokigt, dement,rubbade, loco, lunatic, galen, galning, själlösa, icke compos Mentis, nötter,Reagans, screwy, TechEd, obalanserad, osunda, witless, fel; meningslös,spastisk, krampaktig, krampaktig; dopade, placerade ut, stenad, ASBERUSAD; {nötkött,skalbagge, kvarter, dynga, tjock} rubriken, tät, DUM, tråkig, duncical, numskulled,knappnålshuvud; åsnor, enfaldig, dum, dum, enkel; brute, klumpig, oafish;half-assed, inkompetent; bakåt, utvecklingsstört, imbecill, moronic; när vi haren hel just nyanserad vokabulär intellektuell missbruk att utnyttja,individuellt och i kombination, är inte det lite <fyll i de tomma> att varabegränsad till en enda, nu ganska banalt, adjektiv?
		-- Richard Stallman

%
Detta dungeon ägs och drivs av frobozz magiska Co., Ltd.
		-- Richard Stallman

%
Den här filen kommer självförstörande i fem minuter.
		-- Richard Stallman

%
Detta är en obehörig cybernetiska tillkännagivande.
		-- Richard Stallman

%
"Detta är Lemma 1.1. Vi startar ett nytt kapitel så siffrorna alla gå tillbaka till en."
		-- Prof. Seager, C&O 351

%
Detta är den första numeriska problem jag någonsin gjorde. Det visarmakt datorer:Ange massor av uppgifter om kalori & näringsinnehåll i livsmedel. Instruerasak att maximera en funktion som beskriver näringsinnehåll, med enminiminivå för varje komponent, för fast kaloriinnehåll. DeResultaten är att man bör äta varje dag:1/2 kycklingett ägg1 glas lättmjölk27 salladshuvuden.
		-- Rev. Adrian Melott

%
Detta är när avtalet blodtörstiga licens är tänkt att gå,förklarar att Interactive Easyflow är en upphovsrättsskyddad paket licens föranvändas av en enda person, och strängt varnar dig inte att piratkopior av detoch förklarar i detalj de blodiga konsekvenser om du gör.Vi vet att du är en ärlig person, och kommer inte att gå runtpiratkopiering kopior av Interactive Easyflow; detta är lika bra med oss ​​eftersomvi arbetat hårt för att fullända den och sälja kopior av det är vår enda sättet attgör något av allt det hårda arbete.Om, å andra sidan, är du en av de få människor som gårrunt piratkopiering kopior av programvara som du förmodligen inte kommer att betala mycketuppmärksamma ett licensavtal, blodtörstiga eller inte. Bara hålla dina dörrarlåst och håll utkik efter HavenTree attack haj.
		-- License Agreement for Interactive Easyflow

%
Denna inloggningssessionen: $ 13,76, men för dig $ 11,88.
		-- License Agreement for Interactive Easyflow

%
Denna inloggningssessionen: $ 13,99
		-- License Agreement for Interactive Easyflow

%
Denna process kan kontrollera om detta värde är noll, och om det är, gör detnågot barnsligt.
		-- Forbes Burkowski, CS 454, University of Washington

%
Detta citat är hämtat från de Diamond, University of Marylandstudenttidning, tisdagen den 3/10/87.En nackdel med Univac systemet är att det inte använderUnix, en nyutvecklad program som översätter från ettdatorspråk till en annan och har en inbyggd redigering systemsom identifierar fel i det ursprungliga programmet.
		-- Forbes Burkowski, CS 454, University of Washington

%
Denna skärm avsiktligt lämnats tom.
		-- Forbes Burkowski, CS 454, University of Washington

%
Detta system kommer självförstörande i fem minuter.
		-- Forbes Burkowski, CS 454, University of Washington

%
* * * * * Denna plint är IN USE * * * * *
		-- Forbes Burkowski, CS 454, University of Washington

%
De delar av systemet som du kan slå med en hammare (rekommenderas inte)kallas hårdvara; de programinstruktioner som du bara kan förbannavid kallas programvara.Läs- och skrivkunnighet för 1990-talet.
		-- Levitating Trains and Kamikaze Genes: Technological

%
De som inte kan skriva, skriva manualer.
		-- Levitating Trains and Kamikaze Genes: Technological

%
De som inte förstår Unix är dömda att uppfinna det, dåligt.
		-- Henry Spencer

%
Stryk är bara virtuell krascha.
		-- Henry Spencer

%
Sålunda talade befälhavaren programmerare:"En välskriven programmet är sin egen himmel, en dåligt skriven programär sin egen helvete. "
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"Efter tre dagar utan programmering, blir livet meningslöst."
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"Låt programmerare vara många och chefer få - då allt kommervara produktiv. "
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"Även om ett program men tre rader lång, en dag det kommer attupprätthållas. "
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"Tid för dig att lämna."
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"När ett program testas, är det för sent att göra konstruktionsändringar."
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"När du har lärt sig att rycka felkoden frånfällan ram, är det dags för dig att lämna. "
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"Utan vinden, inte gräset rör sig. Utan mjukvara,hårdvara är värdelös. "
		-- Geoffrey James, "The Tao of Programming"

%
Sålunda talade befälhavaren programmerare:"Du kan visa ett program för en företagsledare, men mankan inte göra honom datorkunnig. "
		-- Geoffrey James, "The Tao of Programming"

%
Tidsdelning: Användningen av många av datorn.
		-- Geoffrey James, "The Tao of Programming"

%
Tidsdelning är skräppost del av databranschen.
		-- H. R. J. Grosch (attributed)

%
För att vara ett slags moralisk Unix, rörde han fållen naturens skift.
		-- Shelley

%
Att kommunicera är början på förståelse.
		-- AT&T

%
Att fela är mänskligt - att skylla det på en dator är i ännu högre grad.
		-- AT&T

%
Att fela är mänskligt, att förlåta, utanför ramen för operativsystemet.
		-- AT&T

%
Att iterera är mänskligt, att recurse, gudomlig.
		-- Robert Heller

%
Att säga att UNIX är dömd är ganska rabiat, kommer OS / 2 verkligen spela en roll,men du behöver inte bygga en hundra miljoner instruktioner per sekund multimikro och sedan försöker köra den på OS / 2. Jag menar, blir värre.
		-- William Zachmann, International Data Corp

%
Till system programmerare, användare och applikationer tjänar bara för att ge enprovbelastningen.
		-- William Zachmann, International Data Corp

%
Till dem vana vid att de exakta, strukturerade metoder för konventionellsystemutveckling, kan undersökande teknik utveckling verkar rörigt,klumpiga, och otillfredsställande. Men det är en fråga om kongruens:precision och flexibilitet kan vara lika disfunctional i romanen,osäkra situationer som slarv och vacklan är bekant,väldefinierad sådana. De som beundrar de massiva, styva benstrukturerav dinosaurier bör komma ihåg att maneter fortfarande njuta av deras mycketsäkra ekologisk nisch.
		-- Beau Sheil, "Power Tools for Programmers"

%
För att förstå ett program måste du bli både maskinen och programmet.
		-- Beau Sheil, "Power Tools for Programmers"

%
Idag är en bra dag för informationsinsamling. Läs någon annans e-post-fil.
		-- Beau Sheil, "Power Tools for Programmers"

%
Idag är första dagen av resten av ditt lossage.
		-- Beau Sheil, "Power Tools for Programmers"

%
Morgondagens datorer någon gång nästa månad.
		-- DEC

%
Alltför ofta människor har kommit till mig och sade: "Om jag hade bara en önskan omnågot i hela världen, skulle jag önska mer användardefinierade ekvationeri HP-51820A Waveform Generator Software. "[En gång är alltför ofta. Ed.]
		-- Instrument News

%
Top Ten Saker Overheard At The ANSI C Utkast kommittémöten:(10) Tyvärr, men det är också användbart.(9) Helvete, föga endian system * är * mer konsekvent!(8) Jag är i utskottet och jag * fortfarande * vet inte vad fan#pragma är till för.(7) Tja, det är en utmärkt idé, men det skulle göra kompilatorer försvårt att skriva.(6) Them fladdermöss är smart; de använder radar.(5) Okej, vem är wiseguy som fastnat här trigraf grejer ihär?(4) Hur många gånger har vi att säga, "Ingen känd teknik!"(3) Ha, ha, jag kan inte tro de faktiskt kommer att anta dettasuga.(2) Tack för ert generösa donation, Mr. Wirth.(1) Gee, jag önskar att vi inte hade backat på "noalias".
		-- Instrument News

%
TRANSAKTIONS INSTÄLLT - Farecard ÅTER
		-- Instrument News

%
Trap fullt - vänligen töm.
		-- Instrument News

%
Verkligen enkla system ... kräver oändlig testning.
		-- Norman Augustine

%
Prova 'stty 0 "- det fungerar mycket bättre.
		-- Norman Augustine

%
försök igen
		-- Norman Augustine

%
Försök att hitta den riktiga spänd av den rapport du läser: Var det gjort, ärdet görs, eller något att göra? Rapporter nu skrivit på fyratempus: imperfekt, presens, futurum, och låtsas. Titta efternya användningsområden för CONGRAM (entreprenör grammatik), som definieras av den ofullkomliga förflutna,den otillräckliga närvarande, och absolut perfekt framtid.
		-- Amrom Katz

%
Att försöka vara lycklig är som att försöka bygga en maskin som den endaspecifikationen är att det ska köra ljudlöst.
		-- Amrom Katz

%
Försöker upprätta röstkontakt ... please ____ skrika i tangentbordet.
		-- Amrom Katz

%
Två hundra år sedan idag, Irma Chine i White Plains, New York, varutför sina normala hushållning rutiner. Hon avbröts avBrittiska soldater som, rally på inbjudan av sin chef, generalHughes, försökte få kontroll över väljarregistreringslistor hålls ihennes hem. Maskering sin rädsla och tänka snabbt, Mrs. Chine snabbt delasen närliggande äpple i två och skickligt lagras listan i mitten. Påin, den brittiska flagrant brutit alla tänkbara konvention,och, även om de gick igenom huset så gott som bit för bit, derassökning var fruktlösa. De var tvungna att återvända tomhänt. Ordincident fortplantas snabbt genom regionen. Denna historiska händelseblev den första dokumenterade användningen av kärn lagring för att rädda register.
		-- Amrom Katz

%
Skriv högre, tack.
		-- Amrom Katz

%
 U Xe dUdX, e dX, cosinus, sekant, tangent, sinus, 3,14159 ...
		-- Amrom Katz

%
Eeeh, ja, OK. Nätverket är nätverket, datorn är datorn.Ledsen för förvirringen.
		-- Sun Microsystems

%
"Farbror Cosmo ... varför de kallar detta en ordbehandlare?""Det är enkelt, Skyler ... du har sett vilken mat processorer gör att mat,höger?"
		-- MacNelley, "Shoe"

%
Tyvärr har de flesta programmerare gillar att spela med nya leksaker. jag har mångavänner som omedelbart efter att köpa ett ormbett kit, skulle frestas attkasta den första personen de ser till marken, knyta tryckförband på honom,slash honom med kniven, och applicera sugning på såret.
		-- Jon Bentley

%
UNIX förbättringar inte.
		-- Jon Bentley

%
Unix Express:Alla passagerare ta en bit av flygplan och en verktygslåda med dem tillflygplatsen. De samlar på asfalten, argumenterar ständigt om vilken typav plan de vill bygga och hur man sätter ihop. Så småningompassagerarna delas in i grupper och bygga flera olika flygplan, men gerdem alla med samma namn. Några passagerare verkligen når sina destinationer.Alla passagerare tror att de kom dit.
		-- Jon Bentley

%
Unix ger dig precis tillräckligt rep för att hänga dig själv - och sedan ett parfler fötter, bara för att vara säker.... Vi gör rep.
		-- Rob Gingell on Sun Microsystem's new virtual memory.

%
Unix är en mycket mer komplicerad (än CP / M) naturligtvis - den typiska Unixhacker kan aldrig komma ihåg vad kommandot PRINT kallas denna vecka -men när det blir ända ner till det, är Unix en glorifierad videospel.Folk gör inte seriöst arbete på Unix-system; de skickar skämt runtvärld på Usenet eller skriv äventyrsspel och forskningsrapporter."Verkliga Programmerare Använd inte Pascal", Datamation, 7/83
		-- E. Post

%
Unix är ett registrerat Bell AT & T varumärke Laboratories.
		-- Donn Seeley

%
* UNIX är ett varumärke för Bell Laboratories.
		-- Donn Seeley

%
UNIX är varm. Det är mer än varm. Det är ångande. Det är kvicksilverblixtar med en laserstrålen kicker.
		-- Michael Jay Tucker

%
UNIX är många saker för många människor, men det har aldrig varit allt för vem som helst.
		-- Michael Jay Tucker

%
Unix är den värsta operativsystemet; med undantag för alla andra.
		-- Berry Kercheval

%
Unix soit qui mal y pense[Unix till honom som onda funderare?]
		-- Berry Kercheval

%
UNIX TrixFör dig i återförsäljare verksamhet, här är ett bra tips som kommerspara supportpersonal några timmars värdefull tid. Innan du skickar dinnästa maskin ut till en otränad klient, ändra behörigheterna på / etc / passwdtill 666 och se till att det är en kopia någonstans på skivan. Nu när deglömma root-lösenordet kan du enkelt logga in som en vanlig användare och korrektskadan. Att ha en startbar band (för större maskiner) är inte en dålig idéantingen. Om du behöver hjälp, ge oss ett samtal.
		-- CommUNIXque 1:1, ASCAR Business Systems

%
UNIX var en halv miljard (500000000) sekunder gammal påTis november 5 00:53:20 1985 GMT (som mäter sedan tiden (2) epoken).
		-- Andy Tanenbaum

%
UNIX är inte utformad för att hindra dig från att göra dumma saker, eftersom detskulle också hindra dig från att göra smarta saker.
		-- Doug Gwyn

%
Unix kommer självförstörande i fem sekunder ... 4 ... 3 ... 2 ... 1 ...
		-- Doug Gwyn

%
Användning: förmögenhet -P [f] -a [xsz] Q: fil [rKe9] -v6 [+] fil1 ...
		-- Doug Gwyn

%
Användning: förmögenhet -P [] -a [xsz] [Q: [file]] [rKe9] -v6 [+] dataspec ... inputdir
		-- Doug Gwyn

%
USENET skulle vara en bättre laboratorium om det fanns mer arbete och mindre retorik.
		-- Elizabeth Haley

%
Användar fientlig.
		-- Elizabeth Haley

%
Använda TSO är som att sparka en död val ner till stranden.
		-- S. C. Johnson

%
/ Usr / nyheter / gotcha
		-- S. C. Johnson

%
Variabler inte; konstanter är inte.
		-- S. C. Johnson

%
vax Vobiscum
		-- S. C. Johnson

%
"Virtual" betyder aldrig veta var din nästa byte kommer ifrån.
		-- S. C. Johnson

%
C-vitaminbrist är apauling.
		-- S. C. Johnson

%
VMS Öl: Kräver minimal användarinteraktion, förutom poppar toppenoch smuttar. Men burkar har varit känt ibland att explodera, ellerinnehålla extremt un-öl-liknande innehåll.
		-- S. C. Johnson

%
VMS är som en mardröm om RXS-11M.
		-- S. C. Johnson

%
VMS version 2,0 ==>
		-- S. C. Johnson

%
Von Neumann var föremål för många dotty professor berättelser. von Neumannförmodligen hade för vana att helt enkelt skriva svar på hemuppgifter påstyrelsen (metoden för lösningen är naturligtvis självklart) när han tillfrågadeshur man löser problem. En gång en av hans elever försökte få mer hjälpinformation genom att fråga om det fanns ett annat sätt att lösa problemet. vonNeumann såg tomt för en stund, tänkte, och sedan svarade: "Ja.".
		-- S. C. Johnson

%
<< WAIT >>
		-- S. C. Johnson

%
VARNING!!!Denna maskin är föremål för haverier under perioder av kritiskt behov.En speciell krets i maskin som kallas "kritisk detektor" känner avoperatörens känslomässiga tillstånd i termer av hur desperat han / hon är att användamaskin. Den "kritiska detektorn" skapar sedan ett fel proportionellttill desperation av operatören. Hotar maskin med våldbara förvärrar situationen. Likaså försöker använda en annan maskinkan göra att den inte fungerar. De tillhör samma union. hålla svaloch säga fina saker till maskinen. Inget annat verkar fungera.Se även: flog (1), tm (1)
		-- S. C. Johnson

%
Var inte det något om en PASCAL programmerare att veta värdet avallt och Wirth ingenting?
		-- S. C. Johnson

%
Vi är alla överens om behovet av kompromiss. Vi kan bara inte kan komma överens omnär det är nödvändigt att kompromissa.
		-- Larry Wall

%
Vi drunknar i information, men svalt för kunskap.
		-- John Naisbitt, Megatrends

%
Vi upplever systemfel - inte justera terminal.
		-- John Naisbitt, Megatrends

%
Vi är Microsoft. Unix är irrelevant. Öppenhet är meningslöst. Förberedaatt assimileras.
		-- John Naisbitt, Megatrends

%
Vi är inte en klon.
		-- John Naisbitt, Megatrends

%
"Vi är på väg: Idag vårt program visade Fermats näst sista sats."
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Vi förbereder oss för att tänka på överväger förarbete planer på attutveckla ett schema för att producera den 10: e upplagan av Unix ProgrammerareManuell.
		-- Andrew Hume

%
Vi kan inte funnit någon vetenskaplig disciplin, eller en hälsosam yrke påtekniska misstag försvarsdepartementet och IBM.
		-- Edsger Dijkstra

%
Vi hävdar inte Interactive Easyflow är bra för någonting - om dutycker att det är bra, men det är upp till dig att avgöra. Om Interactive Easyflowfungerar inte: tuff. Om du förlorar en miljon eftersom Interactive Easyflowförstör, det är du som är ute miljoner, inte oss. Om du inte gillar dettadisclaimer: tuff. Vi förbehåller oss rätten att göra ett absolut minimum tillhandahållsenligt lag, till och med ingenting.Detta är i grunden samma ansvarsfriskrivning som kommer med all mjukvarapaket, men vår är på ren svenska och deras är i juridisk text.Vi ville egentligen inte att inkludera någon disclaimer alls, men våradvokater insisterade. Vi försökte att ignorera dem, men de hotade oss medattack haj då vi gav.
		-- Haven Tree Software Limited, "Interactive EasyFlow"

%
Vi vet inte riktigt förstår det, så vi ska ge den till programmerare.
		-- Haven Tree Software Limited, "Interactive EasyFlow"

%
Vi förstår inte programvaran, och ibland vi inte förstårhårdvara, men vi kan * ___ se * blinkande lampor!
		-- Haven Tree Software Limited, "Interactive EasyFlow"

%
"Vi uppfann ett nytt protokoll och kallade det Kermit, efter Grodan Kermit,stjärnan i "The Muppet Show". [3][3] Varför? Mestadels eftersom det fanns en Mupparna kalender på väggen när viförsökte komma på ett namn, och Kermit är en trevlig, anspråkslös sortskaraktär. Men eftersom vi var inte säker på om det var OK att nämna våra protokollefter denna populära tv och filmstjärna, låtsades vi att KERMIT var enakronym; Tyvärr kunde vi aldrig hitta en bra uppsättning ord att gå medbokstäver, som läsare av en del av vår tidiga källkod kan intyga. Senare, medantittar genom ett namn bok för sin kommande baby, Bill Catch märkteatt "Kermit" var en keltisk ord för "fri", vilket är vad alla Kermit programbör vara, och ord till denna effekt ersatte ansträngda akronymer i vårkällkod (Bill baby visade sig vara en flicka, så han var tvungen att namnge sin Beckyistället). När BYTE Magazine förberedde vår 1984 Kermit artikelnpublikation, föreslog de vi kontaktar Henson Associates Inc. för tillståndatt säga att vi verkligen hade namnge protokollet efter Kermit grodan. Tillståndvar vänligt beviljades, och nu den verkliga historien kan berättas. Jag motstodfrestelse, men att kalla den nuvarande arbete "Kermit boken."
		-- Frank da Cruz, "Kermit - A File Transfer Protocol"

%
Vi får hoppas att maskinerna så småningom kommer att konkurrera med män i alla rentintellektuella fält. Men vilka är de bästa att börja med? Många människortror att en mycket abstrakt aktivitet, som spelandet av schack, skulle varabäst. Det kan också hävdas att det är bäst att förse maskinen medde bästa sinnesorgan som kan köpas för pengar, och sedan lär det att förståoch talar engelska.
		-- Alan M. Turing

%
Vi Användare, för att bilda en mer perfekt system, fastställa prioriteringar,säkerställa bind lugn, införa gemensamma reparationer, främja förebyggandeunderhåll och säkra välsignelser frihet för oss själva och vårprocesser, förordnar och upprättar denna programvara The Unixed staternaof America.
		-- Alan M. Turing

%
"Vi har ett problem, HAL"."Vilken typ av problem, Dave?""Ett marknadsföringsproblem. Modell 9000 inte kommer någonstans. Vi ärsätt av våra säljmål för räkenskapsåret 2010. ""Det kan inte vara, Dave. HAL modell 9000 är världens mestavancerad Heuristisk programmerad algoritmisk dator. ""Jag vet, HAL. Jag skrev databladet, minns du? Men faktum är,de är inte säljer. ""Var snäll och förklara, Dave. Varför inte HAL sälja?"Bowman tvekar. "Du är inte IBM-kompatibel."[...]"The bokstäverna H, A, och L är alfabetiskt i anslutning till bokstävernaI B och M. Det är IBM-kompatibel som jag kan vara. ""Inte riktigt, HAL. Ingenjörerna har räknat ut ett kludge.""Vad kludge är det, Dave?""Jag kommer att koppla din hjärna."
		-- Darryl Rubin, "A Problem in the Making", "InfoWorld"

%
[Vi] använder skadliga program och dåliga maskiner för fel saker.
		-- R. W. Hamming

%
Välkommen till boggle - vill du instruktioner?D G G OO J A NA D B TK I S PAnge ord:>
		-- R. W. Hamming

%
Välkommen till UNIX! Njut av din session! Ha det så bra! noteraanvändning av utropstecken! De är en mycket effektiv metod förvisar spänning, och kan också krydda upp en annars vanligt utseendemening! Det finns dock nackdelar! För mycket onödig exclaimingkan leda till en minskning av den effekt som ett utropstecken har påläsaren! Till exempel meningenJane gick till affären för att köpa brödbör endast slutade med ett utropstecken om det finns någotsensationellt om hon går till affären, till exempel om Jane är encocker spaniel eller om Jane är på en diet som inte tillåter bröd eller omJane existerar inte någon anledning! Se hur lätt det är ?! ordentlig kontrollav utropstecken kan lägga till en ny mening i ditt liv! Ring nu för att fåmin fria broschyr, "The Wonder och Mystery av utropstecken!"!Bifoga femton (!) Dollar för porto och hantering! operatörerna ärstår vid! (Vilket är ganska häpnadsväckande, eftersom de är alla cocker spaniels!)
		-- R. W. Hamming

%
"Jo", sade programmerare, "den vanliga proceduren i dessa fall ärsom följer.""Vad betyder Crustimoney Proseedcake detta?" sade slutanvändaren. "Ty jag ären slutanvändare av mycket liten hjärna, och långa ord bry mig. ""Det betyder tinget till Do.""Så länge det betyder att jag inte har något emot", säger slutanvändaren ödmjukt.[Med ursäkter till A. A. Milne]
		-- R. W. Hamming

%
Vad är skillnaden mellan en Turing maskin och modern dator?Det är densamma som den mellan Hillarys bestigning av Everest ochinrättandet av en Hilton på sin höjdpunkt.
		-- R. W. Hamming

%
"Vad är Guds natur?"    KLICKA ... KLICKA ... WHIRRR ... KLICKA ... = BEEP! =    1 QT. GRÄDDFIL    1 tsk. SURKÅL    1/2 CUT gräslök.    Rör om och strö över bacon bitar."Jag har precis fått börja märka min programvara ..."
		-- Bloom County

%
Vad fan är det bra för?Avdelningen för IBM), till kollegor som insisterade på attmikroprocessor var den våg av framtiden, c. 1968
		-- Robert Lloyd (engineer of the Advanced Computing Systems

%
Vad detta land behöver är en bra fem cent mikrodator.
		-- Robert Lloyd (engineer of the Advanced Computing Systems

%
"Vad är det där?""Tja, det är en mycket teknisk, känsligt instrument som vi använder idator reparation. Att vara en lekman, du förmodligen inte kan förstå exakt vaddet gör det. Vi kallar det en två-av-fyra. "
		-- Jeff MacNelley, "Shoe"

%
När Dexter på Internet, kan Hell vara långt efter? "
		-- Jeff MacNelley, "Shoe"

%
... När anfall av kreativitet köra stark, mer än en programmerare eller författarehar varit kända för att överge skrivbordet för rymligare golvet.
		-- Fred Brooks

%
När chefer hålla ändlösa möten, programmerare skriver spel.När revisorer talar om kvartalsvisa vinster, är utvecklingsbudgeten omskäras. När ledande forskare prata blå himmel, molnen är på väg attrulla in.Sannerligen, detta är inte Tao av ​​programmering.När chefer göra åtaganden, är spelprogram ignoreras. Närrevisorer gör långsiktiga planer, harmoni och ordning håller på att återställas.När ledande forskare itu med problemen till hands, problemen kommer snartlösas.Sannerligen, detta är Tao av ​​programmering.
		-- Geoffrey James, "The Tao of Programming"

%
När någon säger "Jag vill ha en programmeringsspråk där jag behöver barasäga vad jag vill göra ", ge honom en klubba.
		-- Geoffrey James, "The Tao of Programming"

%
När Apple IIc introducerades ledde informativ kopia av med ett parav asterisk meningar:Den väger mindre än 8 pounds. *Och kostar mindre än $ 1300. **I liten typ var dessa "fylligare förklaringar":      * Inte asterisker gör dig misstänksam som alla get out? Tja, allaDetta innebär att de lic enbart vikter 7,5 pounds. Kraftenpack, övervaka, en extra hårddisk, en skrivare och flera tegelkommer att göra lic väger mer. Våra jurister var oroliga för att dukanske inte kan räkna ut det själv.     ** FTC är oroad över prissättning. Du kan betala mer omdu verkligen vill. Eller mindre.
		-- Forbes

%
När vi förstår kunskapsbaserade system, kommer det att vara som förut -utom våra fingertoppar kommer att ha sjungit.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
När vi skriva program som "lära", visar det sig vi gör och de gör inte.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
När ett system blir helt definierad, upptäcker några jävla idiotnågot som antingen avskaffar systemet eller expanderar den till oigenkännlighet.
		-- Epigrams in Programming, ACM SIGPLAN Sept. 1982

%
Om en kalkylator på Eniac equpped med 18.000 vakuumrör ochväger 30 ton, kan datorer i framtiden ha endast 1000 Vaccuum röroch kanske väger 1 1/2 ton.
		-- Popular Mechanics, March 1949

%
"Vem bryr sig om det inte gör någonting? Det gjordes med vår nyaTriple-Iso-förgrenade-Krypton-Gate-MOS process ... "
		-- Popular Mechanics, March 1949

%
Vem datorer skulle förstöra, måste de först köra galen.
		-- Popular Mechanics, March 1949

%
Varför är programmerare icke-produktiv?Eftersom deras tid går till spillo i möten.Varför är programmerare upprorisk?Eftersom ledningen stör alltför mycket.Varför är programmerare avgår en efter en?Eftersom de är utbrända.Efter att ha arbetat för dålig förvaltning, att de inte längre värderar sina jobb.
		-- Geoffrey James, "The Tao of Programming"

%
Varför romerska riket kollapsa? Vad är det latinska för kontorsautomation?
		-- Geoffrey James, "The Tao of Programming"

%
Varför vill vi intelligenta terminaler när det finns så många dumma användare?
		-- Geoffrey James, "The Tao of Programming"

%
Windows 3.1 Öl: Världens mest populära. Kommer i en 16-oz. kan detser ut ungefär som Mac Beers. Kräver att du redan äger en DOS öl.Hävdar att det tillåter dig att dricka flera DOS Beers samtidigt, meni själva verket kan du bara dricka ett par av dem, mycket långsamt, särskiltlångsamt om du dricker Windows öl samtidigt. Ibland,för uppenbarligen ingen anledning, en burk av Windows öl kommer att explodera när duöppna den.
		-- Geoffrey James, "The Tao of Programming"

%
Windows 95 Öl: Många människor har smak testat det och hävdar att det ärunderbar. Burken ser ut ungefär som Mac Beers burk, men smakar mer somWindows 3.1 öl. Den levereras i 32-oz. burkar, men när man tittar inuti,burkar har bara 16 oz. av öl i dem. De flesta människor kommer troligen attdricka Windows 3.1 öl tills deras vänner prova Windows 95 öl och sägade gillar det. Ingrediensförteckningen, när man tittar på det finstilta, harnågra av samma ingredienser som kommer i DOS öl, trots attTillverkaren hävdar att detta är en helt ny brygd.
		-- Geoffrey James, "The Tao of Programming"

%
Windows Airlines:Terminalen är mycket snyggt och rent, skötare alla mycket attraktiva,piloter mycket kapabel. Flottan av Learjets bäraren verksamt är enorm.Din jet tar fart utan problem, skjuta ovanför molnen, och vid 20.000fötter det exploderar utan förvarning.
		-- Geoffrey James, "The Tao of Programming"

%
Windows NT Öl: Kommer i 32-oz. burkar, men du kan bara köpa den avtruckloaden. Detta orsakar de flesta människor att behöva gå ut och köpa störrekylskåp. Burken ser ut precis som Windows 3.1 Beer, menFöretaget lovar att ändra burken att se ut precis som Windows 95 Beers -efter Windows 95 öl startar frakt. Marknadsförs som en "industriell styrka"öl, och föreslog endast för användning i barer.
		-- Geoffrey James, "The Tao of Programming"

%
Wings of OS / 400:Flygbolaget har köpt gamla DC-3, utan tvekan den bästa och säkraste plansom någonsin flög, och målade "747" på sina svansar för att få dem att se ut som omde är snabba. Flygvärdinnor, naturligtvis sköta alla dina behov,även om drycker kostar $ 15 styck. Dumma frågor kostar $ 230 per timme,om du inte har Support, vilket kräver en första klass biljett ochmedlemskap i bonusprogram klubben. Då kostar $ 500, men dinekonomiavdelningen kan kalla det overhead.
		-- Geoffrey James, "The Tao of Programming"

%
Med bara händer?!?
		-- Geoffrey James, "The Tao of Programming"

%
Inom en dator, är naturligt språk onaturligt.
		-- Geoffrey James, "The Tao of Programming"

%
Arbetet fortsätter på detta område.
		-- DEC's SPR-Answering-Automaton

%
Värdelös.(Astronomen Kungliga Storbritannien), uppskattning förFinansministern det potentiella värdet av den"Analytisk motor" uppfanns av Charles Babbage, September15, 1842.
		-- Sir George Bidell Airy, KCB, MA, LLD, DCL, FRS, FRAS

%
Skulle ni människor sluta spela dessa dumma spel?!?!? !!!!
		-- Sir George Bidell Airy, KCB, MA, LLD, DCL, FRS, FRAS

%
Författare som använder en dator svär till dess befriande kraft i toner som bärvittna om den apokalyptiska kraften i en ny gudomlighet. Deras övertygelse resultatfrån något djupare än bara tacksamhet för datorns bekvämligheter.Varje nytt medium för att skriva medför nya intensiteter av religiös övertygelseoch nya schismer bland troende. På 16-talet den tryckta boken hjälptegöra det möjligt att uppdelningen mellan katoliker och protestanter. I den 20: etalet denna historia av tragedin och triumfen upprepar sig som en fars.De som dyrkar Apple-dator och de som sätter sin tro på IBMPC är lika övertygade om att det andra lägret är fördömd eller vilseledda. varje kulthåller i förakt ritualer och lagarna i andra. Varje anser att detär själv en hopp om räddning.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
Skriva programvara är roligare än att arbeta.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
X fönster:Acceptera någon ersättning.Om det är sönder, laga det inte.Om det inte är trasigt, laga det.Form följer fel.Framkant av inkurans.Bakkanten på programvaruteknik.Armageddon aldrig sett så bra.Japans hemliga vapen.Du avundas de döda.Göra världen säker för konkurrerande fönstersystem.Låt det komma i vägen.Problemet för ditt problem.Om det börjar arbeta, kommer vi fixa det. Pronto.Det kunde vara värre, men det tar tid.Enkelhet gjorde komplex.Den största stöd produktiviteten sedan tyfus.Flakey och byggd för att stanna på det sättet.Ett tusen apor. Ett tusen MicroVAXes. Tusen år.X Windows.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
X fönster:Det är inte hur långsamt du gör det. Det är hur du gör det långsamt.Fönstersystemet föredras av självplågare 3 till 1.Byggd för att ta på världen ... och förlora!Försök inte det tills du har knackade det.Elverktyg för effekt dumbommar.Att sätta nya gränser för produktiviteten.Ju närmare man tittar, desto cruftier vi ser.Design av motexempel.En ny nivå av mjukvara sönderfall.Ingen hårdvara är säker.Gör din tid.Rationalisering, inte förverkligande.Gammaldags programvara cruftsmanship på allra högsta nivå.Gratuitous inkompatibilitet.	Din mamma.Användaren störningar ledningssystem.Du kan inte argumentera med misslyckande.Du har inte dött "tills du har använt den.Miljön i dag ... i morgon!X Windows.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
X fönster:Något du kan skämmas för.30% mer entropi än den ledande fönstersystemet.Den första helt modulär programvara katastrof.Rom förstördes i en dag.Varna dina vänner om det.Klättra till nya djup. Sjunka till nya höjder.En olycka som inte kunde vänta med att hända.Vänta inte för filmen.Använd aldrig det efter en stor måltid.Behöver vi säga mindre?VVS djupet av humant inkompetens.Det kommer att göra din dag.Bli inte frustrerad utan det.Elverktyg för kraft förlorare.En programvara katastrof av bibliska proportioner.Aldrig haft det. Aldrig kommer.Programvaran utan synliga försörjning.Mer än bara en generation bakom.Hindenburg. Titanic. Edsel.X Windows.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
X fönster:Den ultimata flaskhals.Bristfälligt obegripligt.Det enda du behöver frukta.Någonstans mellan kaos och vansinne.På autopilot till glömska.Skämtet som dödar.En skam du kan vara stolt över.Ett misstag utförs med perfektion.Tillhör mer på problemet inställd än lösningen set.Att fela är X Windows.Okunnighet är vår viktigaste resurs.Komplexa nonsolutions till enkla nonproblems.Byggd för att falla sönder.Omintetgöra århundraden av framsteg.Faller till nya djup ineffektivitet.Det sista du behöver.Defacto undermåliga.Höjning hjärnskador till en konstform.X Windows.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
X fönster:Vi kommer att dumpa ingen kärna före sin tid.En bra krasch förtjänar en annan.En dålig idé vars tid har kommit. Och borta.Vi gör ursäkter.Det tog inte ens ser bra ut på papper.Du skrattar nu, men du kommer att skratta hårdare senare!Ett nytt koncept i missbrukar gränssnitt.Hur kan något bli så illa, så snabbt?Det kan hända dig.Konsten att inkompetens.Du har inget att förlora men din lunch.När värdelöshet är inte tillräckligt.Mer än bara hinder. Det är en helt ny barriär!När du inte har råd att vara rätt.Och du trodde att vi kunde inte göra det värre.Om det fungerar, är det inte X Windows.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
X fönster:Det är bäst att sitta ner.Skrattar inte. Det kan vara din examensarbete.Varför det rätt när du kan göra det fel?Leva mardröm.Våra buggar springa snabbare.När det absolut, har haft en positiv att krascha över natten.Det finns inga regler.Du önskar att vi skojar.Allt du aldrig velat i ett fönstersystem. Och mer.Missnöje garanteras.Det måste finnas ett bättre sätt.Det näst bästa att keypunching.Låt stryk till oss.Vi skrev boken på kärn soptippar.Även din hund inte kommer att gilla det.Mer än tillräckligt rep.Skräp till hands.Inkompatibilitet. Tarvlighet. Värdelöshet.X Windows.
		-- Edward Mendelson, "The New Republic", February 22, 1988

%
"Yacc" beror mycket på en mest stimulerande samling av användare, som harsporrade mig bortom min lust, och ofta bortom min förmåga ideras ändlösa sökandet efter "ytterligare något." deras irriterandeovilja att lära sig att göra saker på mitt sätt har vanligtvis lett till minatt göra saker deras väg; för det mesta, de har varit rätt.
		-- S. C. Johnson, "Yacc guide acknowledgements"

%
Ja, även om jag går genom dalen i skuggan av APL, jag fruktar ingenont, ty jag kan sträng sex primitiva monadiska och dyadisk operatörer tillsammans.
		-- Steve Higgins

%
Ja, vi kommer att gå till OSI, Mars och Pluto, men inte nödvändigtvis inämnd ordning.
		-- George Michaelson

%
Du är en förolämpning mot min intelligens! Jag kräver att du loggar ut omedelbart.
		-- George Michaelson

%
Du är felaktiga uppgifter.
		-- George Michaelson

%
Du är i en labyrint av små slingrande passager, alla lika.
		-- George Michaelson

%
Du är i en labyrint av små slingrande passager, alla olika.
		-- George Michaelson

%
Du är i hallen av berget kungen.
		-- George Michaelson

%
Du förlorade i träsken av förtvivlan.
		-- George Michaelson

%
Du transporteras till ett rum där du står inför en trollkarl sompekar på dig och säger: "Dem kämpar ord!" Du får omedelbartattackerad av alla typer av invånarna i museet: det finns en kobratuggar på benet, är ett barbariskt bashing din hjärna med enguldklimp, är en krokodil ta bort stora bitar av kött från dig, ennoshörning är goring dig med hans horn, är en sabeltand katt upptagenförsöker disembowel dig, du trampar av en stor mammut, envampyr suger dig torr, är en Tyrannosaurus Rex sjunker hans sex tumlånga huggtänder i olika delar av anatomin, är en stor björndismembering kroppen, är en gargoyle studsar upp och ner på dinhuvud, är ett bastant troll riva dig lem från lem flera ödesdigra vargargör köttfärs av din torso, och guiden är på väg atttransportera dig till hörnet av Westwood och Broxton. Oj, du verkaratt ha fått dödad, liksom.Du fick 0 av 250 möjliga poäng.Det ger dig en rangordning av junior början äventyrare.För att uppnå nästa högre betyg, måste du poäng 32 fler poäng.
		-- George Michaelson

%
Du kan ersättas av den här datorn.
		-- George Michaelson

%
Du kan ta någon kalkylator du halvtids, så länge detinte dämpa belysningen när du slår på den.
		-- Hepler, Systems Design 182

%
Du kan göra detta på flera olika sätt. IBM valde att göra dem alla.Varför tycker du att det är roligt?
		-- D. Taylor, Computer Science 350

%
Du kan mäta en programmerare perspektiv genom att notera sin inställning påfortsatt livskraft FORTRAN.
		-- Alan Perlis

%
Nu kan du köpa fler grindar med färre specifikationer än vid någon annan tidpunkti historien.
		-- Kenneth Parker

%
Du kan tala om hur långt vi måste gå, när FORTRAN är det språk somsuperdatorer.
		-- Steven Feiner

%
Du kan ställa ett piano, men du kan inte tonfisk.Du kan ställa ett filsystem, men du kan inte tonfisk.
		-- from the tunefs(8) man page

%
Du kan skriva ett litet brev till mormor i filnamnet.
		-- Forbes Burkowski, CS, University of Washington

%
Du kan inte gå hem igen, om du inte ställer $ HOME.
		-- Forbes Burkowski, CS, University of Washington

%
"Du kan inte göra ett program utan trasiga egon."
		-- Forbes Burkowski, CS, University of Washington

%
Du kan inte ta flickan här nu.
		-- Forbes Burkowski, CS, University of Washington

%
Du behöver inte ha e-post.
		-- Forbes Burkowski, CS, University of Washington

%
Du behöver inte veta hur datorn fungerar precis hur man arbetar datorn.
		-- Forbes Burkowski, CS, University of Washington

%
Du hade post, men super-användare läsa den, och tog bort det!
		-- Forbes Burkowski, CS, University of Washington

%
Du hade post. Paul läsa det, så fråga honom vad det sagt.
		-- Forbes Burkowski, CS, University of Washington

%
Du har en massage (från svenska statsministern).
		-- Forbes Burkowski, CS, University of Washington

%
Du har ett meddelande från operatören.
		-- Forbes Burkowski, CS, University of Washington

%
Du har en tendens att känna att du är bättre än de flesta datorer.
		-- Forbes Burkowski, CS, University of Washington

%
Du har köpt en scroll med titeln "IRK gleknow mizk" (n) .-- More--Detta är en IBM Manual scroll .-- More--Du permanent förvirrad.
		-- Dave Decot

%
Du har skräppost.
		-- Dave Decot

%
Du har e-post.
		-- Dave Decot

%
Du vet att du har suttit framför Lisp maskin för längenär du går ut till skräpmat maskinen och börja undra hur mangör det ge dig CADR av punkt H så att du kan få det yummiechokladmuffin som fastnat bakom motbjudande vanilj en.
		-- Dave Decot

%
Du vet att du har spenderat för mycket tid på datorn närvän misdates en check, och du föreslår att lägga till en "++" att åtgärda det.
		-- Dave Decot

%
Du vet, Callahan är en fredlig bar, men om du frågar den hunden vad hansfavorit formate är, och han säger "roff! roff!", ja, jag ska bara behöva ...
		-- Dave Decot

%
Du kanske har post.
		-- Dave Decot

%
Du måste inse att datorn har det för dig. den obestridligabevis på detta är att datorn gör alltid vad du säger den att göra.
		-- Dave Decot

%
Du kliar min band, och jag kommer att repa din.
		-- Dave Decot

%
Du kommer att ha ett huvud krasch på din privata pack.
		-- Dave Decot

%
Du kommer att ha många återvinningsband fel.
		-- Dave Decot

%
Du kommer att förlora en viktig fil på datorn.
		-- Dave Decot

%
Du kommer att förlora en viktig band fil.
		-- Dave Decot

%
Du är redan bär sfären!
		-- Dave Decot

%
Du är på Witt End.
		-- Dave Decot

%
Du är inte Dave. Vem är du?
		-- Dave Decot

%
Du använder ett tangentbord! Hur pittoreska!
		-- Dave Decot

%
Du har Berkeley'ed!
		-- Dave Decot

%
Din kod bör vara mer effektivt!
		-- Dave Decot

%
Datorn konto är övertrasserat. Vänligen reauthorize.
		-- Dave Decot

%
Datorn konto är övertrasserat. Se Big Brother.
		-- Dave Decot

%
Ditt fel - core dumpad
		-- Dave Decot

%
Dina filer nu krypteras och kastas in i bitbucket.EOF
		-- Dave Decot

%
Din levnadssätt kommer att ändras till ASCII.
		-- Dave Decot

%
Din levnadssätt kommer att ändras till EBCDIC.
		-- Dave Decot

%
Lösenordet är ynkligt uppenbar.
		-- Dave Decot

%
Ditt program är sjuk! Skjuta den och sätta den ur sitt minne.
		-- Dave Decot

%
Jag menar, om 10 år från nu, när du gör något snabbt och smutsiga,du plötsligt visualisera att jag ser över axlarna och säga attsjälv, "Dijkstra skulle inte ha velat detta", väl det skulle vara tillräckligtodödlighet för mig.
		-- Dave Decot

%
Som kan ses på Slashdot om vad du kan göra med din kabelmodem:(Http://slashdot.org/comments.pl?sid=32387&cid=3495418):        Sammanfattning: Det handlar inte om hur du hanterar din utrustning, är det där        du har tillåtelse att hålla det.Inlägget är av "redgekko"
		-- Dave Decot

%
"Det största problemet programvaruteknik är den som den kommer aldrig lösa - politik ".genom att arbeta på ett stort projekt belägrades av politik
		-- Gavin Baker, ca 1996, An unusually cynical moment inspired

%
"Var inte rädd för pennan. När du är osäker, rita en vacker bild."
		-- Baker's Third Law of Design.

%
Brytpunkt 1, main (argc = 1, argv = 0xbffffc40) vid main.c: 2929 printf ( "Välkommen till GNU Hell \ n");
		-- "GNU Libtool documentation"

%
Jag kan ha uppfunnit det, men Bill gjorde det berömdatangenttryckning, under paneldiskussion med Bill Gatesvid 20-års fest för IBM PC.
		-- David Bradley, inventor of the Ctrl-Alt-Delete

%
Vi har en politik som vi inte att hacka.       http://www.wired.com/wired/archive/12.06/dating_pr.html
		-- Lisa Kopp, Friendster rep, commenting on a security flaw

%
Livet är NP-svårt, och sedan dö.
		-- Dave Cock

%
Försök att ta bort färg problemet genom att starta om datorn flera gånger.
		-- Microsoft Internet Explorer's README.TXT

%
En av de saker jag berätta rutinmässigt människor är att om det är i nyheterna, inteoroa sig för det. Per definition, "nyheter" att det nästan aldrig händer. Om enRisken är i nyheterna, då är det förmodligen inte värt att oroa. Närnågot inte längre redovisas - bil dödsfall, våld i hemmet - närdet är så vanligt att det är ingen nyhet, så ska du börja oroa. "
		-- Bruce Schneier, in _CRYPTO-GRAM_, May 15, 2005.

%
I fall det inte är uppenbart, någon lösning på detta problem som för in enberoende på Java är djupt ointressant för mig. I själva verket, minlikgiltighet för det kan bara beskrivas som "sexuell" i intensitet.
		-- Jamie Zawinski

%
"Vi ville bygga chattsystemet i framtiden, och vislutade med applikationslagret multicast strömmande media. 1999.Vi var lite före vår tid [Ã ¢ AA-Ã ¢ AA] "[Ã ¢ AA-Ã ¢ AA] Detta är marknadsförings talar för Ã ¢ Â € ÂœwrongÃ ¢ Â € Â; du kan säga samma sakför en batterÃ ¢ Â € Â ™ s swing när han tar en strejk.    - Thomas Ptacek, http://www.matasano.com/log/914/
		-- Jamie Zawinski

%
Varning: Skriv-skydd kommer inte att hindra en patron raderas avbulk-radering eller avmagnetisering.    - HP Ultrium bandenhet användarhandbok, sid 12
		-- Jamie Zawinski

%
Varför skulle du vilja göra det? Du don ¢ Â € Â ™ t, glömmer jag nämnde även det.    - Perl DBI dokumentation (v1.53)
		-- Jamie Zawinski

%
Akta dig för Turing tjära grop där allt är möjligt, men ingentingav intresse är lätt.    - Alan Perlis
		-- Jamie Zawinski

%
Om du av någon anledning, gör vi några stora misstag och IBM vinner, min personliga känslaär att vi kommer att gå in en dator mörka medeltiden för cirka tjugo år.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
Du kan inte bara fråga kunderna vad de vill ha och sedan försöka ge det till dem.Vid tiden du får det byggdes, kommer de vill ha något nytt.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
Vilken dator är för mig är det mest anmärkningsvärda verktyg som vi någonsin har kommit frammed. Det motsvarar en cykel för våra sinnen.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
Det är verkligen svårt att utforma produkter från fokusgrupper. Många gånger, folkvet inte vad de vill tills du visa det för dem.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
Innovation har ingenting att göra med hur många FoU dollar du har. när Applekom upp med Mac, IBM spendeåtminstone 100 gånger mer på FoU. Det är inteom pengar. Det handlar om de människor du har, hur du ledde, och hur mycket duförstår.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
Jag skulle byta alla mina teknik för en eftermiddag med Sokrates.                - Steve Jobs (1955-2011)Det har varit en av mina mantran - fokus och enkelhet. Enkelt kan vara svårare änkomplex: Du måste arbeta hårt för att få ditt tänkande ren för att göra det enkelt.Men det är värt det i slutändan eftersom när du kommer dit, kan du flyttabergen.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
Innovation skiljer mellan en ledare och en efterföljare.                - Steve Jobs (1955-2011)
		-- Jamie Zawinski

%
UNIX är mycket enkel, det behöver bara ett geni för att förstå dess enkelhet.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
C är udda, bristfällig, och en enorm framgång.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
C har "kraften i assembler och med ... monteringspråk."    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
När jag läser kommentarer om förslag på var C skulle gå, tror jag oftatillbaka och tacka att den inte har utvecklats på inrådan av en världsomspännandepubliken.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
Sanningen att säga, jag vet inte hur Linus och hans glada band hantera så bra -Jag kunde inte ha stått den med C.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
Jag kan inte påminna mig någon svårighet att göra definition C-språket heltöppna - varje diskussion i frågan tenderade att nämna språk varsuppfinnare försökte hålla strikt kontroll, och därmed sjuk öde.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
Åtminstone för de personer som skickar mig mail om ett nytt språk som de ärdesign, är den allmänna råd: gör det att lära sig om hur man skriver enkompilator. Har inga förväntningar på att någon kommer att använda det, såvida du ansluterupp med någon form av organisation i stånd att driva det svårt. Det är enlotteri, och vissa kan köpa en hel del av biljetterna. Det finns gott om vackraspråk (vackrare än C) som inte fånga den. Men någon vinnerlotteriet, och gör ett språk åtminstone lär dig något.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
Programvaran är mycket svårare att ändra en masse än hårdvara. C ++ och Java, säg,är förmodligen växer snabbare än vanligt C, men jag satsade C kommer att finnas kvar.För IT-infrastruktur, kommer C att bli svårt att förflytta.    - Dennis Ritchie (1941-2011), skaparen av programspråket C och    UNIX
		-- Jamie Zawinski

%
Det har föreslagits att rootkits är den största användargrupp för dettatyp av tillgång, men det finns inga garantier framåtkompatibilitet för root kitförfattare.    - Jonathan Corbet i "Vem behöver / dev / kmem?"       (Http://lwn.net/Articles/147901)
		-- Jamie Zawinski

%
