(1) Kontors anställda dagligen sopa golv, damma avmöbler, hyllor och montrar.(2) Varje dag fyller lampor, rena skorstenar, och trimma vekar.Tvätta fönstren gång i veckan.(3) Varje kontorist kommer att medföra en hink med vatten och en ventilationsluckor avkol för dagens verksamhet.(4) Gör din pennor noggrant. Du kanske skära spetsar till dinindividuell smak.(5) Detta kontor öppnas klockan 07:00 och stänger vid 08:00 utompå sabbaten, på vilken dag vi kommer att förbli stängd. Varjeanställd förväntas tillbringa sabbaten genom att närvarakyrka och bidra frikostigt till orsaken till Herren.Works, 1872
		-- "Office Worker's Guide", New England Carriage

%
(6) män anställda kommer att ges ledigt varje vecka för att uppvaktaändamål, eller två kvällar i veckan om de går regelbundet i kyrkan.(7) Efter en anställd har tillbringat sina tretton timmars arbete ikontor, skulle han tillbringa den återstående tiden läsa Bibelnoch andra goda böcker.(8) Varje anställd bör lägga undan från varje betala paket en ansenligsumman av sina resultat för hans fördel under sina sjunkande år,så att han inte kommer att bli en börda för samhället eller hans betters.(9) En anställd som röker spanska cigarrer, använder alkoholhaltig drycki någon form, frekventerar biljardbord och offentliga hallar, eller blirrakat i en frisör butik, kommer att ge mig goda skäl att misstänkahans värd, avsikter, integritet och ärlighet.(10) Den anställde som har utfört sitt arbete troget ochutan fel under fem år, kommer att få en ökning avfem cent per dag i hans lön, som ger vinster frånföretag tillåter det.
		-- "Office Worker's Guide", New England Carriage Works, 1872

%
En bank är en plats där de ger du ett paraply i vackert väder ochbe om det tillbaka när det börjar regna.
		-- Robert Frost

%
En chef utan humor är som ett jobb som är inget kul.
		-- Robert Frost

%
En budget är bara en metod för att oroa innan du spenderar pengar, samtsom efteråt.
		-- Robert Frost

%
En affärsman är en hybrid av en dansare och en miniräknare.
		-- Paul Valery

%
Ett utskott är en grupp som håller minuter och förlorar timmar.
		-- Milton Berle

%
Ett utskott är en livsform med sex eller fler ben och ingen hjärna.
		-- Lazarus Long, "Time Enough For Love"

%
En kommitté slår rot och växer, den blommar, wilts och dör, spridning avutsäde från vilka andra utskott kommer att blomma.
		-- Parkinson

%
En kommun är där människor går samman för att dela deras brist på rikedom.
		-- R. Stallman

%
Ett företag är känd av män det håller.
		-- R. Stallman

%
En konsult är en person som lånar din klocka, berättar vilken tid detär, fickor klockan, och skickar en faktura för det.
		-- R. Stallman

%
En fortsatt flöde av papper är tillräcklig för att fortsätta pappersflödet.
		-- Dyer

%
En ko är en helt automatiserad mjölktillverkningsmaskin. Den är inkapsladi ogarvade skinn och monterade på fyra vertikala, rörliga stöden, en vidvarje hörn. Den främre änden av maskinen, eller inmatning, innehåller den skärandeoch slipmekanism, som utnyttjar en unik återkopplingsanordning. Även här ärstrålkastarna, luftintag och avgas en stötfångare och en mistlur.Baktill på maskinen bär den mjölk utmatningsutrustning somsamt en inbyggd ominspelade och insekts repeller. Den centrala deleninrymmer en hydro kemisk-omvandlingsenheten. I korthet består detta av fyrajäsning och lagringstankar seriekopplade genom ett intrikat nätverkflexibel VVS. Denna enhet innehåller också den centrala värmeanläggningenkomplett med automatiska temperaturkontroll, pumpstation och huvudventilationssystem. Apparaten avfalls ligger på baksidan avdenna mittsektion.Kor är tillgängliga fullt monterade i ett sortiment av storlekar ochfärger. Produktionen varierar från 2 till 20 ton mjölk per år. Ikorthet de viktigaste yttre synliga detaljer i kon är: två åskådare, tvåfnask, fyra stander-överdelar, fyra hängare-Downers, och en swishy-wishy.
		-- Dyer

%
En matnings försäljare är på väg till en gård. Som han kör längs på fyrtioen magisterexamen, han ser ut sin bil fönstret och ser en trebent kyckling igångtillsammans med honom, hålla jämna steg med sin bil. Han är förvånad över att en kyckling ärkörs vid fyrtio en magisterexamen Så han hastigheter upp till fyrtiofem, femtio, då sextioen magisterexamen Kycklingen håller rätt upp med honom hela vägen, sedan plötsligtlyfter och försvinner i fjärran.Mannen drar in på gården och säger till bonden, "Du vet,den märkligaste just hänt mig; Jag körde längs vid åtminstonesextio miles i timmen och en kyckling passerade mig som om jag stod stilla! ""Ja", bonden svarar, "det kyckling var vårt. Du ser, det finnsmig, och det finns Ma, och det är vår son Billy. När vi hade kyckling förmiddag, skulle vi alla ha en trumpinne, så vi skulle behöva döda två kycklingar.Så vi bestämde att försöka föda upp en trebent kyckling så var och en av oss kundehar en trumpinne. ""Hur smakar de?" sade bonden."Vet inte", svarade bonden. "Vi har inte kunnat fångaen ännu. "
		-- Dyer

%
En frilans är en som får betalt av ordet - per styck eller kanske.
		-- Robert Benchley

%
En bra handledare kan trampa på tårna utan stöka din glans.
		-- Robert Benchley

%
Ett holdingbolag är en sak där du lämnar en medbrottsling varorna medanpolisen söker dig.
		-- Robert Benchley

%
En man är bekant vid företaget som han anordnar.
		-- Ambrose Bierce

%
Ett möte är ett evenemang där minuterna hålls och timmar förlorade.
		-- Ambrose Bierce

%
En promemoria skrivs inte informera läsaren, utan för att skydda författaren.
		-- Dean Acheson

%
En motion att ajournera är alltid i ordning.
		-- Dean Acheson

%
En mus är en elefant som byggs av japanerna.
		-- Dean Acheson

%
En ny leverans av runda tuits har kommit och är tillgängliga från Mary.Någon som har skjutit upp arbetet tills de fick en rundatuit nuhar ingen ursäkt för ytterligare förhalning.
		-- Dean Acheson

%
En rock butik så småningom stängas; de tog för mycket för granit.
		-- Dean Acheson

%
... Något som heter Etik, vars natur var förvirrande men om du hade det duvar en hög klass fastighetsmäklare och om du hade inte du var en shyster, en piker ochen fly-by-night. Dessa dygder väckt förtroende och möjligt för dig att hanteraStörre Propositions. Men de inte innebära att du skulle vara opraktisktoch vägrar att ta dubbelt så mycket för ett hus om en köpare var en sådan idiotatt han inte tvinga dig ner på det begärda priset.
		-- Sinclair Lewis, "Babbitt"

%
En resande försäljare körde förbi en gård när han såg en gris med treträben utför en magnifik serie backflips och hjula.Förbryllad, körde han upp till gården, där han hittade en gammal bondesitter på gården tittar grisen."Det är ganska en gris du har där, sir", sa försäljaren."Visst är, son," bonden svarade. "Varför, för två år sedan, min dottervar simma i sjön och stötte huvudet och förbannat nära drunknade, men attgris simmade ut och drog henne tillbaka till stranden. ""Fantastiskt!" försäljaren utropade."Och det är inte det enda. I höstas var jag Cuttin trä upp pånorra fyrtio när ett träd föll på mig. Nålas mig till marken, gjorde det.Det gris köra upp och vickade under trädet och lyfte den av mig.Räddade mitt liv.""Fantastiskt! Försäljaren sa. Men säg mig, hur kommer grisen hartre träben? "Bonden stirrade på nykomlingen i förvåning. "Mister, när dufick en amazin "gris som att du inte äta honom alla på en gång."
		-- Sinclair Lewis, "Babbitt"

%
Ett muntligt avtal är inte värt papperet det är skrivet på.
		-- Samuel Goldwyn

%
Om den tid som vi tror att vi kan gå ihop, någon flyttar ändarna.
		-- Herbert Hoover

%
Enligt en färsk och ovetenskaplig nationell undersökning, leende är någotalla bör göra minst 6 gånger per dag. I ett försök att ökanationella genomsnittet (USA rankas på tredje plats bland världens stormakter iler), har Xerox instruerat all personal att vara glad, sprudlande, ochviktigast av allt, att le. Xerox medarbetare är överens om, och även känna starktatt de inte bara kan träffas utan att överträffa det nationella genomsnittet ... utom förTubby Ackerman. Men eftersom Tubby gör en sådan bra jobb med racing runtparkeringsplatser med en stor fjäril netto hämta flytande IC-chips, Xeroxbeslutade att ge honom en paus. Om du ser Tubby på en parkeringsplats han kan haen fåraktigt flin. Det är där uttrycket "Service med en någotsheepish flin "kommer från.
		-- Herbert Hoover

%
Enligt alla de senaste rapporterna, fanns det ingen sanning i någon avtidigare rapporter.
		-- Herbert Hoover

%
Reklam är en värdefull ekonomisk faktor eftersom det är den billigastesätt att sälja varor, särskilt om varorna är värdelösa.
		-- Sinclair Lewis

%
Reklam är rasslande en pinne i en matavfall hink.
		-- George Orwell

%
Reklam kan beskrivas som vetenskapen om att arrestera mänskligaintelligens tillräckligt länge för att få pengar från det.
		-- George Orwell

%
När allt är sagt och gjort, är en fan av mycket mer sagt än gjort.
		-- George Orwell

%
Efter någon lön höjning, kommer du att ha mindre pengar i slutet avmånad än vad du gjorde innan.
		-- George Orwell

%
Allt jag begär är en chans att bevisa att pengar kan inte göra mig lycklig.
		-- George Orwell

%
Alla de stora företagen depreciera sina ägodelar, och du kan också,förutsatt att du använder dem i affärssyfte. Till exempel, om du prenumererarWall Street Journal, en företagsrelaterade tidningen kan du dra avkostnaden för ditt hus, eftersom det i ord US Supreme Court ChiefJustice Warren Burger i ett landmärke 1979 skattebeslut: "Var annars är dukommer att läsa tidningen? Utanför? Vad händer om det regnar? "
		-- Dave Barry, "Sweating Out Taxes"

%
Allt detta big deal om ekonomisk brottslighet - vad är det för fel med vit kragebrottslighet? Som trivs med sitt jobb idag? Du? Mig? Vem som helst? Den enda tillfredsställandedel av alla jobb är kaffepaus, lunch timme och avsluta tid. För flera år sedanDet var åtminstone hopp om förbättring - eventuella främjande - merviktiga jobb framöver. När du kan säljas myten om att du kan göraVD för företaget du nästan aldrig stjäla frimärken. men ingentror han kommer att bli president längre. Ju fler människor byter jobbju mer de inser att det finns ett direkt samband mellan att arbeta fören levande och total bedövande tristess. Så varför inte ta hämnd? Du är intekommer att hitta mig knackar en kille eftersom han kuddar ett utgiftskonto och hanshem pappers bär företagets emblem. Ta bort brott från den vitaTjänsteman och du kommer att beröva honom hans sista resten av jobbet intresse.
		-- J. Feiffer

%
Allt detta mygel runt, varför, är det inte för pengarna, är det för skojs skull.Pengar är precis som vi räkna poäng.
		-- Henry Tyroon

%
Alla säkerhets- och garantiklausuler blir ogiltigt vid betalning av fakturan.
		-- Henry Tyroon

%
Amerika fungerar mindre, när du säger "Union ja!"
		-- Henry Tyroon

%
Amerikanska näringslivet länge sedan gav upp kräver att blivande anställdavara ärlig och hårt arbetande. Det har till och med slutat hoppas för anställda som ärutbildade nog att de kan skilja mellan män rummet ochdamernas rum utan lite bilder på dörrarna.
		-- Dave Barry, "Urine Trouble, Mister"

%
Ett kontor parti är inte, som ibland tänkt verkställande direktörenschans att kyssa te-flicka. Det är te-flickans chans att kyssaVD (dock bisarra ambitionen detta kan verka till någonsom har sett VD ansikte på).
		-- Katherine Whitehorn, "Roundabout"

%
Vem som helst kan göra någon mängd arbete under förutsättning att det är inte det arbete han är tänktatt göra just nu.
		-- Robert Benchley

%
Vem som helst kan hålla rodret när havet är lugnt.
		-- Publius Syrus

%
Vem som helst kan göra en omelett med ägg. Tricket är att göra en med ingen.
		-- Publius Syrus

%
Något gratis är värt vad du betalar för det.
		-- Publius Syrus

%
Allt märkt "NY" och / eller "förbättrade" är inte. Etiketten innebärpriset gick upp. Etiketten "ALLA NYA", "HELT NY", eller "Stora nya"innebär att priset gick upp.
		-- Publius Syrus

%
"Åtminstone de är ___________ ERFARNA incompetents"
		-- Publius Syrus

%
Vid dessa priser, jag förlorar pengar - men jag gör det upp i volym.
		-- Peter G. Alaquon

%
På jobbet är omvänt proportionell mot den av en personantal pennor som personen bär.
		-- Peter G. Alaquon

%
Vara social. Tala med personen bredvid dig i arbetslöshetlinjen i morgon.
		-- Peter G. Alaquon

%
Förts sistone?
		-- Peter G. Alaquon

%
... Innan jag kunde komma till någon slutsats slog det mig att mitt taleller min tystnad, faktiskt några åtgärder till mig, skulle vara en ren meningslöshet. Vadgjorde det roll vad någon visste eller ignoreras? Vad betydde det som varchef? Man får ibland en sådan blixt av insikt. Det viktigaste idenna affär låg djupt under ytan, bortom räckhåll, och bortom minmakt inblandning.
		-- Joseph Conrad

%
Mellan 1950 och 1952, en uttråkad meterolog, stationerad norr om HudsonBay, lämnade ett monument som varken regeringen eller tid kan utrota.Med hjälp av en bulldozer övergiven av flygvapnet, tillbringade han två år ochstor möda trycka stenblock i ett enda ord.Det kan ses från 10.000 fot, silhuett mot snön.Regeringstjänstemän utbytte PM full av omskrivningar (ingen latinmotsvarande existerar) men misslyckades med att uttrycka ett anslag räkningen förförstörelse av detta röse, skulle det inte varna pressen och generabåde parlamentet och Party.Det står i dag, ett monument till mänskliga anden. Om liv existerar på andraplaneter, kan detta vara det första meddelandet som mottagits från oss.
		-- The Realist, November, 1964.

%
Akta dig för alla företag som kräver nya kläder, och inte hellreen ny bärare av kläder.
		-- Henry David Thoreau

%
Biz är bättre.
		-- Henry David Thoreau

%
Body av Nautilus, Brain av Mattel.
		-- Henry David Thoreau

%
Bullwinkle: Du lämnar just det till min kompis. Han är hjärnan hos kläderna.Allmänt: Vad som gör DU?Bullwinkle: Vad? En verkställande.
		-- Jay Ward

%
Business är ett bra spel - massor av konkurrens och minimum av regler.Du håller poäng med pengar.
		-- Nolan Bushnell, founder of Atari

%
Verksamhet kommer att vara antingen bättre eller sämre.
		-- Calvin Coolidge

%
"Men oroa dig inte, dess för en sak - att mata globala företags tassar."
		-- Calvin Coolidge

%
Men den största Elektrisk Pioneer av dem alla var Thomas Edison, som var enlysande uppfinnare trots att han hade lite formell utbildning ochbodde i New Jersey. Edisons första stora uppfinning i 1877, vargrammofon, som snart kunde hittas i tusentals amerikanska hem, därdet i princip satt fram till 1923, när posten uppfanns. Men Edisonsstörsta bedrift kom 1879, när han uppfann elbolaget.Edison design var en lysande anpassning av enkel elektrisk krets:elbolaget skickar elektricitet genom en kabel till en kund, dåomedelbart får el tillbaka genom en annan tråd, sedan (detta ärden lysande delen) sänder det tillbaka till kunden igen.Detta innebär att en elektrisk företag kan sälja en kund samma partiel tusentals gånger om dagen och aldrig fastna, eftersom mycket fåkunder tar sig tid att undersöka sin el noga. I själva verket denförra året en ny el producerades i USA var 1937;de elbolag har bara åter sälja det sedan dess, vilket ärvarför de har så mycket ledig tid att ansöka om räntehöjningar.
		-- Dave Barry, "What is Electricity?"

%
I mitten av 1880-talet, nästan alla vägar utom de iSyd, var av den nuvarande standarden spårvidd. De sydliga vägarna varfortfarande fem fot mellan skenorna.Det beslutades att ändra spårvidden alla södra vägar till standard,på en dag. Denna anmärkningsvärda arbete utfördes på en söndag majav 1886. I flera veckor i förväg, hade affärer varit upptagen press hjul påaxlar till den nya och smalare spårvidd, att ha ett förråd av rullande materiel somkan köras på det nya spåret så snart som det var klart. Slutligen, den dag som,ett stort antal av gäng av spårlager började arbeta i gryningen. över~~POS=TRUNC allt~~POS=HEADCOMP enjärnväg var lossas, flyttas i tre och en halv inches, och spetsade i sinny position. Genom mörk, tåg från var som helst i USA skulle kunna fungeraöver spåren i söder, och en fritt utbyte av godsvagnar alltvar möjligt.
		-- Robert Henry, "Trains", 1957

%
Genom att arbeta troget åtta timmar om dagen, kan du så småningom få varachef och arbete tolv.
		-- Robert Frost

%
Kan någon komma ihåg när tiderna inte var hårt, och pengar inte knappa?
		-- Robert Frost

%
Kan något vara tråkigare än arbete kvar oavslutade? Ja, arbete aldrig börjat.
		-- Robert Frost

%
Slarvigt planerade projekt tar tre gånger längre tid att slutföra än förväntat.Noggrant planerade projekt ta fyra gånger längre tid att slutföra än förväntat,främst på grund planerarna förväntar sig att deras planering för att minska den tid det tar.
		-- Robert Frost

%
Ordförande i uttråkad.
		-- Robert Frost

%
Kolumn 1 Kolumn 2 Kolumn 30. integrerade 0. ledningen 0. alternativ1. Totalt 1. organisatorisk 1. flexibilitet2. systematiseras 2. övervakas 2. kapacitet3. parallell 3. ömsesidig 3. rörlighet4. funktionell 4. digital programmering 4.5. responsiv 5. logistiskt 5. koncept6. tillval 6. övergångs 6. tids fas7. synkroniserade 7. inkrementell 7. projektion8. kompatibel 8. tredje generationens 8. hårdvara9. balanserad 9. policy 9. beredskapsProceduren är enkel. Tänk på någon tresiffrigt nummer, välj sedanden motsvarande modeord från varje kolumn. Till exempel, nummer 257 producerar"Systematiseras logistiska projektion", en fras som kan släppas inpraktiskt taget alla rapporter med ringen avgörande, kunnig myndighet. "Nejen kommer att ha de mest avlägsna uppfattning om vad du pratar om ", säger Broughton,"Men det viktiga är att de inte är på väg att erkänna det."
		-- Philip Broughton, "How to Win at Wordsmanship"

%
Utskott har blivit så viktigt i dag att underkommittéer måsteutses för att göra jobbet.
		-- Philip Broughton, "How to Win at Wordsmanship"

%
Kompetens, som sanning, skönhet och kontaktlinser, är i ögat avbetraktaren.
		-- Dr. Laurence J. Peter

%
Konkurrenskraftig fury är inte alltid ilska. Det är den sanna missions modoch iver inför möjligheten att ens bästa kanske inte är tillräckligt.
		-- Gene Scott

%
... [Om citattecken] även om vi * ___ gjorde * citat någon i dettaföretag, skulle det förmodligen vara rappakalja.
		-- Thom McLeod

%
"Consequences, Schmonsequences, så länge jag är rik."
		-- "Ali Baba Bunny" [1957, Chuck Jones]

%
Betrakta frimärke: dess användbarhet består i förmågan atthålla sig till en sak tills det blir där.
		-- Josh Billings

%
Konsulter är mystiska människor som frågar ett företag för ett nummer och sedange tillbaka till dem.
		-- Josh Billings

%
Kredit ... är det enda bestående vittnesbörd om människans tilltro till människan.
		-- James Blish

%
Att hantera fel är enkelt:Arbeta hårt för att förbättra.Framgång är också lätt att hantera:Du har löst fel problem.Arbeta hårt för att förbättra.
		-- James Blish

%
Att handskas med problemet med ren personal ackumulation,alla våra undersökningar ... peka på en genomsnittlig ökning på 5,75% per år.
		-- C. N. Parkinson

%
Kära herre:Jag vill bara * ___ en * enarmade manager så jag har aldrig höra "Onandra sidan ", igen.
		-- C. N. Parkinson

%
Kära Mister Språk Person: Vad är syftet med apostrof?Svar: Den apostrof används huvudsakligen i hand märkte små affärer skyltaratt göra läsaren uppmärksam på än ett "S" kommer upp i slutet av ett ord, som i:VI utom inte personlig check'S, eller: EJ ANSVARIG FÖR PUNKT'S.En annan viktig grammatik begrepp att tänka på när du skapar hand bokstävernasmåföretag tecken är att du ska lägga citattecken runt slumpvisord för dekoration, som i "TRY" Hot HUNDS, eller ens försöka "OUR" HOT DOG'S.
		-- Dave Barry, "Tips for Writer's"

%
Trots allt att döma, är din chef en tänkande, känsla, människa.
		-- Dave Barry, "Tips for Writer's"

%
"Tror du vad vi gör är fel?""Det är naturligtvis fel! Det är olagligt!""Jag har aldrig gjort något olagligt innan.""Jag trodde du sa att du var en revisor!"
		-- Dave Barry, "Tips for Writer's"

%
Var inte oersättlig, om du inte kan bytas ut, du kan inte främjas.
		-- Dave Barry, "Tips for Writer's"

%
Stjäl inte; thou'lt aldrig därmed konkurrera framgångsrikt i näringslivet. Fuska.
		-- Ambrose Bierce

%
Säg inte hur hårt du arbetar. Säg mig hur mycket du får gjort.
		-- James J. Ling

%
"Do not tell me jag bränna ljuset i båda ändar - säg mig var attfå mer vax !! "
		-- James J. Ling

%
Drömmar är gratis, men du får dränkts på anslutningstiden.
		-- James J. Ling

%
Borrning efter olja är tråkigt.
		-- James J. Ling

%
Tjäna pengar på din fritid - utpressning dina vänner.
		-- James J. Ling

%
Ernest frågar Frank hur länge han har arbetat för företaget."Ända sedan de hotade att skjuta mig."
		-- James J. Ling

%
Någonsin märker att även de mest trafikerade människor är aldrig för upptagen för att berättahur upptagen de är?
		-- James J. Ling

%
Varje moln har en silverkant; du skulle ha sålt den och köpte titan.
		-- James J. Ling

%
"Varje människa har sitt pris. Mine är $ 3,95."
		-- James J. Ling

%
Varje människa tror Gud är på hans sida. De rika och mäktiga vet att han är.
		-- Jean Anouilh, "The Lark"

%
Varje morgon i Afrika, vaknar en gasell upp. Det vet den måste springa fortareän den snabbaste lejon eller det kommer att dödas. Varje morgon ett lejon vaknar.Det vet den måste springa den långsammaste gasellen eller det kommer att svälta ihjäl.Det spelar ingen roll om du är ett lejon eller en gasell: när solen kommerupp, skulle du bättre vara igång.
		-- Jean Anouilh, "The Lark"

%
"Varje morgon, jag gå upp och titta igenom" Forbes lista överrikaste människorna i Amerika. Om jag inte är där, jag går till jobbet "
		-- Robert Orben

%
Varje framgångsrik person har haft fel, men upprepad underlåtenhet är ingengaranti för eventuell framgång.
		-- Robert Orben

%
Varje ung man bör ha en hobby: att lära sig att hantera pengar ärden bästa.
		-- Jack Hurley

%
Alla men Sam hade anmält sig till ett nytt företag pensionsplan somkallas för en liten anställd bidrag. Företaget betalar allaresten. Tyvärr var 100% anställdas deltagande behövs;annars planen var avstängd. Sam chef och hans arbetskamrater badoch övertalas, men till ingen nytta. Sam sade att planen skulle aldrig löna sig.Slutligen kallas företagets VD Sam in i hans kontor."Sam", sade han, "här är en kopia av den nya pensionsplanen och här ären penna. Jag vill att du ska underteckna papper. Jag är ledsen, men om du inte skriver,du är avskedad. Från och med nu. "Sam tecknat tidningarna omedelbart."Nu", sade presidenten, "skulle du vilja tala om för mig varför dukunde inte har undertecknat tidigare? ""Ja, sir", svarade Sam "ingen förklarade det för mig ganska såklart tidigare. "
		-- Jack Hurley

%
Alla gillar en kidder, men ingen ger honom pengar.
		-- Arthur Miller

%
Alla som kommer in här vill tre saker:(1) De vill det snabbt.(2) De vill ha det bra.(3) De vill ha det billigt.Jag berättar dem att plocka två och ringa mig tillbaka.
		-- sign on the back wall of a small printing company

%
Undantag bekräftar regeln, och förstöra budgeten.
		-- Miller

%
Utdrag ur ett samtal mellan en kundsupport person och enkund som arbetar för en välkänd militär anslutna forskningslaboratorium:Support: "Du är inte vår enda kund, du vet."Kund: "Men vi är en av de få med taktiska kärnvapen."
		-- Miller

%
Executive förmåga beslutar snabbt och få någon annan att göraarbetet.
		-- John G. Pollard

%
Exxons "universum av energi" tenderar att den säregna snarare änhumoristisk ... Efter [en obegriplig film montage om vind och sol ochregn och band gruvor och] två eller tre minuter av mekanisk förvirring, densäten locomote genom en fylld med klockarbets dinosaurier kort tunnel.Dinosaurierna avbildas utan precision och för nära ansiktet."En av de få riktiga nyheter på Epcot är användningen av luktförvärra illusioner. Naturligtvis, ingen vet vad dinosaurierna luktade som,men Exxon har beslutat att de luktade illa."I andra änden av Dino Ditch ... det finns en slutlig, mycket addledmeddelande om att möta challengehood morgon-wise. Jag somnade under denna,men importen verkar vara att dinosaurierna inte har något att göra medenergipolitik och inte heller dig. "
		-- P. J. O'Rourke, "Holidays in Hell"

%
Misslyckande är oftare från brist på energi än brist på kapital.
		-- P. J. O'Rourke, "Holidays in Hell"

%
Snabbt, billigt, bra: plocka två.
		-- P. J. O'Rourke, "Holidays in Hell"

%
Rädsla är den största försäljare.
		-- Robert Klein

%
Känn desillusionerad? Jag har fått några stora nya illusioner, just här!
		-- Robert Klein

%
För varje kille som gör sitt märke, det finns ett halvt dussin väntar på att sudda ut.
		-- Andy Capp

%
Genius är en procent inspiration och nittionio procent svett.
		-- Thomas Alva Edison

%
Genius är tio procent inspiration och femtio vinster procent av kapital.
		-- Thomas Alva Edison

%
Få jobbet gjort är ingen ursäkt för att inte följa reglerna.Naturlig följd:Följa reglerna inte kommer att få jobbet gjort.
		-- Thomas Alva Edison

%
"Med tanke på valet mellan att åstadkomma något och bara ligger runt,Jag skulle snarare ligga runt. Ingen tävling."
		-- Eric Clapton

%
Gud hjälpe dem som inte hjälpa sig själva.
		-- Wilson Mizner

%
Gud hjälper dem som hjälper sig själva.
		-- Benjamin Franklin, "Poor Richard's Almanac"

%
Bra dag för att undvika polisen. Krypa för att arbeta.
		-- Benjamin Franklin, "Poor Richard's Almanac"

%
Bra säljare och bra reparatörer kommer aldrig gå hungrig.
		-- R. E. Schenk

%
Lyckan är ett positivt kassaflöde.
		-- R. E. Schenk

%
Hårt arbete dödade aldrig någon, men varför chansa?
		-- Charlie McCarthy

%
Har du tänkt på att de människor som alltid försöker att berätta`Det finns en tid för arbete och en tid för lek" aldrig hitta tid för lek?
		-- Charlie McCarthy

%
Han har inte fått en förmögenhet; turen har förvärvat honom.
		-- Bion

%
Han som har men fyra och tillbringar fem har inget behov av en plånbok.
		-- Bion

%
Den som är nöjd med sin lott har förmodligen en hel del.
		-- Bion

%
Han som steg på andra för att nå toppen har bra balans.
		-- Bion

%
"Här på telebolaget, vi betjäna alla typer av människor, frånPresidenter och kungar till avskum ... "
		-- Bion

%
"Hej, Sam, vad sägs om ett lån?""Whattaya behöver?""Åh, om $ 500.""Whattaya fick för säkerhet?""Whattaya behöver?""Vad sägs om ett öga?"
		-- Sam Giancana

%
Ohyggligt vanställt av en gammal indisk förbannelse?VI KAN HJÄLPA!Ring (511) 338-0959 för en omedelbar möte.
		-- Sam Giancana

%
Hyra moraliskt handikappade.
		-- Sam Giancana

%
Byggvaruhus är avsedda för gör-det-självare som är villiga attbetala högre priser för att underlätta för att kunna handla timmer,hårdvara och brödrostar alla på ett ställe. Märker jag säga "shop för", sommotsats till "få." Detta är den största nackdelen med hem centra: de äralltid av allt utom konstgjorda julgranar. Hemma centrumanställda har ingen tid att ordna handelsvaror eftersom de är alltför upptagenapplicera litet pris klistermärken på varje objekt - varje bräda, tvättmaskin, spikoch skruva - i hela butiken ...Låt oss säga att en bit i din toalett tank raster, så du tar borttrasiga delen, ta det till hemmet centrum och be en anställd om han har enersättning. Den anställde, som har aldrig sitt liv ens sett insidanav en toalett tank, kommer inbördes vid den trasiga delen i stort sett på samma sättatt en medlem av en primitiv Amazonas djungel stam skulle titta på en elektroniskkalkylator, och sedan säga, "Vi väntar en transport av dessa någon gångi mitten av nästa vecka. "
		-- Dave Barry, "The Taming of the Screw"

%
Ärlighet är för det mesta mindre lönsamt än oärlighet.
		-- Plato

%
Ärlighet lönar sig men det verkar inte betala tillräckligt för att passa vissa människor.
		-- F. M. Hubbard

%
Hotell är trött på att få rippat. Jag checkas in ett hotell och dehade handdukar från mitt hus.
		-- Mark Guido

%
Hur kommer alla kommer så långsamt om det kallas rusningstid?
		-- Mark Guido

%
Hur kommer finansiella rådgivare verkar aldrig vara så rika som dehävdar att de kommer att göra dig?
		-- Mark Guido

%
"Hur många människor arbetar här?""Åh, ungefär hälften."
		-- Mark Guido

%
Mänskliga resurser är mänsklig först och resurser andra.
		-- J. Garbers

%
"Jag är övertygad om att tillverkarna av matt ta bort lukt pulverhar inkluderat inkapslade tid släpptes katt urin i sina produkter.Denna teknik måste vara vad hindrade dess fördelning under min mammasregera. Min matta luktar piss och jag har inte en katt. bättre gåköpa lite mer. "
		-- timw@zeb.USWest.COM

%
Jag är mer uttråkad än du någonsin kan möjligen vara. Gå tillbaka till arbetet.
		-- timw@zeb.USWest.COM

%
Jag tillskriver min framgång till intelligens, mod, beslutsamhet, ärlighet,ambition, och har tillräckligt med pengar för att köpa människor med dessa egenskaper.
		-- timw@zeb.USWest.COM

%
Jag BET det som hände var de upptäckte elden och uppfunnit hjulet påsamma dag. Sedan den natten, brände de hjulet.
		-- Jack Handey, The New Mexican, 1988.

%
Jag kan inte dra en vagn, eller äta torkade havre; Om det är människans arbete jag kommer att göra det.
		-- Jack Handey, The New Mexican, 1988.

%
Jag anser att en ny enhet eller teknik för att ha kulturellt accepterat närDet har använts för att begå ett mord.
		-- M. Gallaher

%
Jag gör det inte för pengarna.
		-- Donald Trump, Art of the Deal

%
Jag har inte någon användning för livvakter, men jag har en specifik användning för tvåvälutbildade auktoriserade revisorer.
		-- Elvis Presley

%
Jag vill inte uppnå odödlighet genom mitt arbete. Jag vill uppnåodödlighet genom att inte dö.
		-- Woody Allen

%
Jag för en kan inte protestera den senaste M.T.A. biljettpris vandra ochåtföljande löften som detta inte på något sätt förbättra servicen. Förtransiteringssystemet, som det nu verkar, har gömt fördelar somkan inte mätas i pengar.Personligen anser jag att det är väl värt 75 cent eller till och med $ 1 tillhar det oantastliga ursäkt när jag är sen till någonting: "Jag kommed tunnelbanan. "Dessa fyra ord har en sådan magi i dem som om Godotbör en dag dyker upp och mumlar dem, någon publik skulle omedelbartförstå sin långa förseningar.
		-- Woody Allen

%
Jag fortsätta att arbeta av samma skäl en höna fortsätter lägga ägg.
		-- H. L. Mencken

%
Jag har de enklaste smaker. Jag är alltid nöjd med det bästa.
		-- Oscar Wilde

%
Jag har sätt att tjäna pengar som du inte vet någonting om.
		-- John D. Rockefeller

%
Jag frågade bara mig själv ... vad skulle John Delorean göra?
		-- Raoul Duke

%
Jag behöver bara tillräckligt för att upptrappade mig tills jag behöver mer.
		-- Bill Hoest

%
Jag gillar arbete; Det fascinerar mig; Jag kan sitta och titta på det i timmar.
		-- Bill Hoest

%
Jag fuskade aldrig en ärlig man, endast rascals. De ville ha något föringenting. Jag gav dem ingenting för något.
		-- Joseph "Yellow Kid" Weil

%
Jag är skyldig allmänheten ingenting.
		-- J. P. Morgan

%
Jag var i detta förtid luftkonditionerade stormarknad och det fanns alladessa gångar och det fanns dessa badmössor du kan köpa som hade dessatyp av fjärde juli putsar på dem som var röd och gul och blå ochJag var inte frestas att köpa en, men jag blev påmind om att jag hade varitundvika stranden.
		-- Lucinda Childs "Einstein On The Beach"

%
Jag var en del av den märkliga ras av människor träffande beskrivits som utgifterderas liv gör saker som de avskyr att tjäna pengar som de inte villköpa saker de inte behöver att imponera på folk de ogillar.
		-- Emile Henry Gauvreay

%
Jag skulle hellre ledas till helvetet än lyckats himlen.
		-- Emile Henry Gauvreay

%
Jag skulle snarare bara tro att det är gjort av små älvor kör runt.
		-- Emile Henry Gauvreay

%
Jag är alltid letar efter en ny idé som kommer att vara mer produktiva än dess kostnad.
		-- David Rockefeller

%
Jag har alla pengar jag någonsin behöver om jag dör av klockan fyra.
		-- Henny Youngman

%
JAG:Det bästa sättet att göra en silke plånbok från en sugga öra är att börjamed en siden sugga. Detsamma gäller pengar.II:Om dagens var hälften så bra som i morgon är tänkt att vara, skulle detförmodligen vara dubbelt så bra som igår var.III:Det finns inga lata veteran lejon jägare.IV:Om du har råd att annonsera, behöver du inte.V:En tiondel av deltagarna producerar mer än en tredjedel av produktionen.En ökning av antalet deltagare minskar bara genomsnittetutgång.
		-- Norman Augustine

%
Om en underordnad ställer en relevant fråga, titta på honom som om han hadeförlorade sina sinnen. När han tittar ner, parafrasera frågan tillbaka på honom.
		-- Norman Augustine

%
Om en sak är värt att göra, är det värt att göra dåligt.
		-- G. K. Chesterton

%
Om en sak är värd att ha, är det värt att fusk för.
		-- W. C. Fields

%
Om allt annat misslyckas, sänka dina normer.
		-- W. C. Fields

%
Om bankirer kan räkna, hur kommer de har åtta fönster och bara fyra rösträknare?
		-- W. C. Fields

%
Om någonsin nöjet att man måste köpas av smärtan av den andra, därbättre vara någon handel. En handel med vilken man får och den andra förlorar är ett bedrägeri.
		-- Dagny Taggart, "Atlas Shrugged"

%
Om Gud inte hade gett oss tejp, skulle det ha varit nödvändigt att uppfinna den.
		-- Dagny Taggart, "Atlas Shrugged"

%
Om jag hade ett gruvschakt, jag tror inte att jag skulle bara överge det. det finnsmåste finnas ett bättre sätt.
		-- Jack Handey, The New Mexican, 1988.

%
Om jag vill ha din åsikt, ska jag be dig att fylla i nödvändiga formen.
		-- Jack Handey, The New Mexican, 1988.

%
Om jag var en dödgrävare eller ens en bödel, det finns vissa människor jag kundearbeta med en stor njutning.
		-- Douglas Jerrold

%
Om det är värt att göra, är det värt att göra för pengarna.
		-- Douglas Jerrold

%
Om pengar inte kan köpa lycka, jag antar att du bara har att hyra den.
		-- Douglas Jerrold

%
Om vi ​​kunde sälja våra erfarenheter för vad de kostar oss, vi skullealla vara miljonärer.
		-- Abigail Van Buren

%
Om vad de har gjort har inte löst problemet, berätta för dem attgöra något annat.
		-- Gerald Weinberg, "The Secrets of Consulting"

%
Om du alltid skjuta nöje du aldrig kommer att få det. Avsluta arbete och spelaför en gångs skull!
		-- Gerald Weinberg, "The Secrets of Consulting"

%
Om du är bra, kommer du att tilldelas allt arbete. Om du är verkligabra, kommer du få ut av det.
		-- Gerald Weinberg, "The Secrets of Consulting"

%
Om du är över 80 år gammal och tillsammans med dina föräldrar, vi kommerlöser in checken.
		-- Gerald Weinberg, "The Secrets of Consulting"

%
Om du fotograferar i 80 du försummar ditt företag;över 80 du försummar din golf.
		-- Walter Hagen

%
Om du inte är rika bör du alltid se bra.
		-- Louis-Ferdinand Celine

%
Om du kan räkna dina pengar, behöver du inte en miljard dollar.
		-- J. Paul Getty

%
Om du inte kan få jobbet gjort under de första 24 timmarna, arbeta nätter.
		-- J. Paul Getty

%
Om du inte kan lära sig att göra det bra, lära sig att njuta av att göra det dåligt.
		-- J. Paul Getty

%
Om du inte behövde jobba så hårt, skulle du ha mer tid att vara deprimerad.
		-- J. Paul Getty

%
Om du gör något rätt en gång, kommer någon ber dig att göra det igen.
		-- J. Paul Getty

%
Om du inte har tid att göra det rätt, där du kommer att hitta tidatt göra det?
		-- J. Paul Getty

%
Om du misslyckas med att planera, planerar att misslyckas.
		-- J. Paul Getty

%
Om du hade bättre verktyg, kan du mer effektivt visa dintotal inkompetens.
		-- J. Paul Getty

%
Om du måste fråga hur mycket det är, kan du inte råd med det.
		-- J. Paul Getty

%
Om du hype något och det lyckas, du är ett geni - det var inte enhype. Om du hype det och det misslyckas, då var det bara en hype.
		-- Neil Bogart

%
Om du säljer diamanter, kan du inte räkna med att ha många kunder.Men en diamant är en diamant, även om det inte finns några kunder.
		-- Swami Prabhupada

%
Om du misstänker att en man, inte anställa honom.
		-- Swami Prabhupada

%
Om du tror att ingen bryr sig om du lever, prova saknas ett par bilbetalningar.
		-- Earl Wilson

%
Om du vill veta vad Gud tänker på pengar, titta bara på de människor han gavdet.
		-- Dorthy Parker

%
Om du vill sätta dig på kartan, publicera din egen karta.
		-- Dorthy Parker

%
Om du vill veta värdet av pengar, gå försöka låna.
		-- Ben Franklin

%
Om du är som de flesta husägare, du är rädd för att många reparationerrunt ditt hem är för svårt att ta itu med. Så när din ugnexploderar, ringer i en så kallad professionell för att fixa det. De"Professionella" anländer i en lastbil med bokstäver på sidorna och avsätter ettstor mängd verktyg och två assistenter som tillbringar större delen av denvecka i källaren handtralla objekt på måfå med tunga skiftnycklar, eftersom "professionella" avkastning och ger dig en faktura för något merpengar än det skulle kosta att driva en framgångsrik kampanj för USASenat.Och det är därför du har beslutat att börja göra saker själv. Dufigur, "Om dessa killar kan fixa min ugn, sedan så kan I. Hur svårt burkdet vara? "	Mycket svårt. De flesta hem projekt är omöjliga, somDärför bör du göra dem själv. Det finns ingen anledning att betala andrafolk att skruva upp saker när du enkelt kan skruva upp dem själv för långtmindre pengar. Den här artikeln kan hjälpa dig.
		-- Dave Barry, "The Taming of the Screw"

%
Viktiga brev som innehåller inga fel kommer att utveckla fel i posten.Motsvarande fel kommer att dyka upp i två exemplar medan Boss läserDet. Vital papper kommer att visa sin vitalitet genom spontant flyttafrån där du lämnade dem till där du inte kan hitta dem.
		-- Dave Barry, "The Taming of the Screw"

%
År 1914 var det första korsord tryckt i en tidning. Deskapare fick $ 4000 ner ... och $ 3000 över.
		-- Dave Barry, "The Taming of the Screw"

%
I konsumtionssamhället finns oundvikligen två typer av slavar:fångarna av missbruk och fångar avund.
		-- Dave Barry, "The Taming of the Screw"

%
I en hierarki varje anställd tenderar att stiga till sin nivå av inkompetens ...i tid varje inlägg tenderar att vara upptagen av en anställd som är inkompetentatt utföra sina uppgifter ... Arbetet utförs av de anställda somhar ännu inte nått sin nivå av inkompetens.
		-- Dr. Laurence J. Peter, "The Peter Principle"

%
Vid atom attack, kommer alla arbets regler tillfälligt.
		-- Dr. Laurence J. Peter, "The Peter Principle"

%
I händelse av skada meddela din chef omedelbart. Han kommer att kyssa den ochgör det bättre.
		-- Dr. Laurence J. Peter, "The Peter Principle"

%
I varje hierarki grädden stiger tills det surnar.
		-- Dr. Laurence J. Peter

%
För att få ett lån måste du först bevisa att du inte behöver det.
		-- Dr. Laurence J. Peter

%
I mitten av ett brett fält är en kruka med guld. 100 fot i norr ståren smart chef. 100 fot i söder står en dum chef. 100 fot tillöst är påskharen, och 100 fot i väst är Santa Claus.Fråga: Vem kommer till kruka med guld först?A: Den dumma manager. Allt annat är myter.
		-- Dr. Laurence J. Peter

%
Innovation är svårt att schemalägga.
		-- Dan Fylstra

%
Insanity är den sista försvar ... Det är svårt att få en återbetalning närförsäljare är sniffa ditt skrev och baying på månen.
		-- Dan Fylstra

%
Är en person som blåser upp banker en econoclast?
		-- Dan Fylstra

%
Det är bättre att ge än att låna ut, och det kostar ungefär samma.
		-- Dan Fylstra

%
Det är bättre att leva rik än att dö rik.
		-- Samuel Johnson

%
Det är bättre att resa förhoppningsvis än att flyga Continental.
		-- Samuel Johnson

%
Det är svårt att sväva med örnarna när du arbetar med kalkoner.
		-- Samuel Johnson

%
Det är absolut nödvändigt när man flyger tränare som du hålla någon tendens tillden levande fantasifulla. För även om det kan momentant verkar varafall är det inte alls sannolikt att kabinen är helt bebos avgråtande barn rökare billiga inhemska cigarrer.
		-- Fran Lebowitz, "Social Studies"

%
Det är omöjligt att njuta av tomgång ordentligt om man har gott omarbete att göra.
		-- Jerome Klapka Jerome

%
Det är mycket svårare att hitta ett jobb än att hålla en.
		-- Jerome Klapka Jerome

%
Det räcker inte att jag skulle lyckas. Andra måste misslyckas.[Också tillskrivas David Merrick. Ed.]Det räcker inte att lyckas. Andra måste misslyckas.[Stora tankar lika? Ed.]
		-- Gore Vidal

%
Det är löjligt att kalla detta en industri. Det här är inte. Detta är råtta äterråtta, hund äter hund. Jag ska döda dem, och jag kommer att döda dem innan dedöda mig. Du pratar om det amerikanska sättet att survival of the fittest.
		-- Ray Kroc, founder of McDonald's

%
Det är en dålig arbetare som skyller sina verktyg.
		-- Ray Kroc, founder of McDonald's

%
Det har varit ett företag gör nöje med dig.
		-- Ray Kroc, founder of McDonald's

%
Det är fantastiskt! Vi har inte sett något liknande i den sista en halvtimme!
		-- Macy's

%
Det är inte så svårt att lyfta sig själv genom dina bootstraps när du är från marken.
		-- Daniel B. Luten

%
Det är väldigt glamoröst att höja miljontals dollar, tills det är dags för denRiskkapitalbolaget att suga dina ögonglober ut.
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Bara för att han är död är inget skäl att avskeda arbete.
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Fortsätt så! Men snälla inte be mig att hjälpa till.
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Håll din chef chef av din chef rygg.
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Håll ögonen på bollen,Axeln till hjulet,Näsan till slipstenen,Fötterna på marken,Ditt huvud på dina axlar.Nu ... försöka få något gjort!
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Påkostade utgifterna kan bli katastrofala. Inte köpa några öser på ett tag.
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Låna ut pengar till en dålig gäldenär och han kommer att hata dig.
		-- Peter Kennedy, chairman of Kraft & Kennedy.

%
Låt mig försäkra er om att för oss här på First National, du är inte bara enantal. Youre två siffror, ett bindestreck, tre fler nummer, en annan streck ochett annat nummer.
		-- James Estes

%
Låt oss organisera denna sak och ta allt det roliga ur det.
		-- James Estes

%
Livet är en hälsosam respekt för moder jord spetsad med girighet.
		-- James Estes

%
Livet är billigt, men tillbehören kan döda dig.
		-- James Estes

%
Leva inom din inkomst, även om du måste låna för att göra det.
		-- Josh Billings

%
Lever på jorden kan vara dyrt, men det finns en årlig gratis resarunt solen
		-- Josh Billings

%
Lo! Män har blivit verktyg för sina verktyg.
		-- Henry David Thoreau

%
Lån avdelningschef: "Det finns inte någon finstilta på dessa.räntor, behöver vi inte det. "
		-- Henry David Thoreau

%
Ensam?Som en förändring?Som ett nytt jobb?Liksom spänning?Gillar att träffa nya och intressanta människor?JUST screw-up EN MER TID !!!!!!!
		-- Henry David Thoreau

%
Titta, vi handla varje dag ute med hustlers, hantera beslutsfattare, shysters,con-män. Det är sättet på vilket företag att komma igång. Det är så härland byggdes.
		-- Hubert Allen

%
Massor av folk förväxla dålig förvaltning med ödet.
		-- Frank Hubbard

%
Kärlek kan skratta åt låssmeder, men han har en djup respekt för pengar påsar.
		-- Sidney Paternoster, "The Folly of the Wise"

%
Lycka, det är då förberedelse och möjlighet möts.
		-- P. E. Trudeau

%
Göra framsteg i arbetet. Fortsätt att låta saker och ting försämras hemma.
		-- P. E. Trudeau

%
Människan är ett djur som gör fynd: inga andra djur gör this--ingen hund byter ben med en annan.
		-- Adam Smith

%
Man måste forma sina verktyg så att de formar honom.
		-- Arthur R. Miller

%
Management: Hur många fötter behöver möss har?Svar: Möss har fyra fötter.M: Utveckla!R: Möss har fem bihang, och fyra av dem är fötter.M: Ingen diskussion av femte bihang!R: Möss har fem bihang; fyra av dem är fötter; en är en svans.M: Vad? Fötter utan ben?R: Möss har fyra ben, fyra fötter och en svans per enhet-mus.M: Förvirrande - är att totalt 9 bihang?R: Möss har fyra ben fot församlingar och en bottenaggregatet per kroppen.M: Inte helt diskutera frågan!R: Varje mus är utrustad med fyra ben och en svans. varje benär utrustad med en fot vid änden motsatt kroppen; svansenär inte utrustad med en fot.M: Beskrivande? Ja. Kraftfull NO!R: Tilldelning av bihang för möss kommer att vara: Fyra fot-ben heter,en svans. Avvikelser från denna policy är inte tillåtet eftersom det skulleutgöra misapportionment knappa bihang tillgångar.M: För auktoritär; kväver kreativitet!R: Möss har fyra fötter; varje fot är fäst på ett litet ben sammanfogadeintegrerat med den övergripande mus strukturella delsystem. Ocksåfäst på mus undersystemet är en tunn svans, icke-funktionella ochprydnadsväxter i naturen.M: För utförlig / vetenskaplig. Svara på frågan!R: Möss har fyra fötter.
		-- Arthur R. Miller

%
Många människor är förtjusta om sitt arbete.
		-- Arthur R. Miller

%
Många människor är förtjusta om ditt arbete.
		-- Arthur R. Miller

%
Många människor skriver PM att berätta de har inget att säga.
		-- Arthur R. Miller

%
Mater Artium necessitas.[Nöden är uppfinningarnas moder].
		-- Arthur R. Miller

%
Föräldrapenning? Nu varje Tom, Dick och Harry blir gravid.
		-- Malcolm Smith

%
Kanske du inte kan köpa lycka, men dessa dagar kan du säkert ladda det.
		-- Malcolm Smith

%
McDonalds - Därför att du är värd det.
		-- Malcolm Smith

%
Män av höga geni när de gör det minst arbete är mest aktiva.
		-- Leonardo da Vinci

%
Män tar endast deras behov i beaktande - aldrig sina förmågor.
		-- Napoleon Bonaparte

%
Män hud skiljer sig från kvinnors hud. Den är vanligen större, ochden har fler ormar tatuerade på den. Dessutom, om du undersöker en kvinnas hudmycket noga, tum för tum, med början på hennes välformade fotleder, sedan försiktigtspåra smal kurva hennes kalvar, sedan flytta upp till henne ...[Redaktörens anmärkning: För att göra plats för nyhetsartiklar om viktiga händelser i världensåsom jordbruk, kommer vi att ta bort de närmaste kvadratfot avkvinnas hud. Tack.]... Tills slutligen två du ligger där, tillbringade, rökning dincigaretter, och plötsligt slår dig: Human hud är faktiskt består avmiljarder små enheter av protoplasma, som kallas "celler"! Och vad som är ännu merintressant, de på utsidan är alla döende! Detta är ett faktum. Dinhud är som en aggressiv modern bolag, där äldre veteranceller, som slutligen har arbetat sig fram till de bästa och erhållna kontormed fin utsikt, ständigt knuffade ut genom fönstret huvudet först,utan så mycket som en pensionsplan, av yngre hotshot celler rör sig upp frånNedan.
		-- Dave Barry, "Saving Face"

%
Mental kraft tenderade att korrumpera och absolut intelligens tenderade attkorrupta absolut, tills offret undvek våld helt iförmån för smarta lösningar på dumma problem.
		-- Piers Anthony

%
Pengar kan inte köpa lycka, men det kan göra dig väldigt bekväm närdu är olycklig.
		-- C. B. Luce

%
Pengar kan inte köpa kärlek, men det förbättrar din förhandlingsposition.
		-- Christopher Marlowe

%
Pengar kan inte köpa kärlek, eller ens vänskap.
		-- Christopher Marlowe

%
Pengar talar inte, det svär.
		-- Bob Dylan

%
Pengar är bättre än fattigdom, om så bara av ekonomiska skäl.
		-- Bob Dylan

%
Pengar är sin egen belöning.
		-- Bob Dylan

%
Pengar är roten till allt ont, och man behöver rötter.
		-- Bob Dylan

%
Pengar är roten till all rikedom.
		-- Bob Dylan

%
Pengar är sanningsenlig. Om en man talar om hans ära, få honom att betala kontant.
		-- Lazarus Long

%
Pengar är inte allt - men det är en lång väg framför vad som kommer härnäst.
		-- Sir Edmond Stockdale

%
Pengar kan köpa vänskap men pengar kan inte köpa kärlek.
		-- Sir Edmond Stockdale

%
Pengar kommer att säga mer i ett ögonblick än de mest vältaliga vännen kan i år.
		-- Sir Edmond Stockdale

%
Moneyliness är bredvid gudaktighet.
		-- Andries van Dam

%
De flesta människor kommer att lyssna på dina orimliga krav, om du ska övervägaderas oacceptabla erbjudande.
		-- Andries van Dam

%
Mundus vult decipi decipiatur ergo.[Världen vill bli lurade, så fuska.]
		-- Xaviera Hollander

%
Min uppfattning om grovbearbetning det är när rumsservice är sent.
		-- Xaviera Hollander

%
Min uppfattning om grovbearbetning det roterande luftkonditioneringen för låg.
		-- Xaviera Hollander

%
Mitt problem ligger i att förena mina brutto vanor med min nettoresultat.Varje människa som har $ 10.000 kvar när han dör är ett misslyckande.
		-- Errol Flynn

%
"Nöden är uppfinningarnas moder" är en dum ordspråk. "Nödvändighetär mor till meningslösa knep "är mycket närmare sanningen.
		-- Alfred North Whitehead

%
Slipsar strypa klart tänkande.
		-- Lin Yutang

%
vädjar aldrig till en mans "bättre natur." Han kanske inte har en.Åberopar sin egennytta ger dig mer inflytande.
		-- Lazarus Long

%
frågar aldrig två frågor i ett affärsbrev. Svaret kommer att diskuteraden du är minst intresserad, och säger ingenting om den andra.
		-- Lazarus Long

%
Aldrig köpa från en rik försäljare.
		-- Goldenstern

%
Aldrig köpa vad du inte vill eftersom det är billigt, kommer det att vara kär för dig.
		-- Thomas Jefferson

%
Ring aldrig en man en dåre. Låna från honom.
		-- Thomas Jefferson

%
Aldrig investera dina pengar i något som äter eller behöver ommålning.
		-- Billy Rose

%
Aldrig hålla jämna steg med de Joneses. Dra ner dem till din nivå.
		-- Quentin Crisp

%
Låt aldrig någon som säger att det inte kan göras avbrott den person som ärgör det.
		-- Quentin Crisp

%
Aldrig säga att du vet en man tills du har delat ett arv med honom.
		-- Quentin Crisp

%
berättar aldrig folk hur man gör saker. Berätta för dem vad de ska göra och de kommeröverraska dig med sin uppfinningsrikedom.
		-- Gen. George S. Patton, Jr.

%
Lita på aldrig någon som säger pengar är inget objekt.
		-- Gen. George S. Patton, Jr.

%
Försök aldrig att lära en gris att sjunga. Det slösar din tid och retar grisen.
		-- Lazarus Long, "Time Enough for Love"

%
NEW YORK-- Kraft Foods, Inc. meddelade idag att dess styrelsedirektörer förkastade enhälligt $ elva miljard maktövertagande bid av PhilipMorris och Co. A Kraft talesman uppgav i en presskonferens atterbjudandet avvisades eftersom det $ 90 per aktie bud inte återspegladesanna värdet av bolaget.Wall Street insiders dock berätta en helt annan historia.Uppenbarligen Kraft styrelse hade alla utom undertecknat övertagandetavtal när de lärt sig av Philip Morris marknadsföringsplaner för en avderas stora Mellanöstern dotterbolag. Till en person, röstade styrelsen attavvisa budet när de upptäckte att tobaksjätten avsedd attomorganisera israeliska Cheddar, Ltd., och namnge det nya bolaget Ost från Nasaret.
		-- Lazarus Long, "Time Enough for Love"

%
Nitwit idéer är för nödsituationer. Du använder dem när du har ingetannat att prova. Om de arbetar, de går i boken. Annars följerBoken, som är i stort sett en samling nitwit idéer som fungerade.
		-- Larry Niven, "The Mote in God's Eye"

%
Ingen kommitté någonsin kunde komma på något så revolutionerande som en kamel -något som är praktiskt möjligt och så perfekt utformad för att fungera effektivt isådana svåra förhållanden.
		-- Laurence J. Peter

%
"Inget jobb för stora, ingen avgift för stor!"
		-- Dr. Peter Venkman, "Ghost-busters"

%
Ingen blir sjuka på onsdagar.
		-- Dr. Peter Venkman, "Ghost-busters"

%
Inga problem är olösligt i alla tänkbara omständigheter.
		-- Dr. Peter Venkman, "Ghost-busters"

%
Inga problem är så formidabel att du inte bara kan gå ifrån det.
		-- C. Schulz

%
Inga problem är så stor att det kan inte vara lämpligt i någonstans.
		-- C. Schulz

%
Inga skidor ta stenar som hyres skidor!
		-- C. Schulz

%
Ingen spotta på bussen!Tack, mgt.
		-- C. Schulz

%
Ingen av våra män är "experter." Vi har mest tyvärr funnit det nödvändigtatt bli av med en man så snart som han tror sig en expert - eftersom ingennågonsin anser sig expert om han verkligen vet sitt jobb. En man som vetjobb ser så mycket mer att göra än vad han har gjort, att han alltid pressarframåt och aldrig ger upp ett ögonblick av tanke till hur bra och hur effektivthan är. Tänker alltid framåt, tänker alltid att försöka göra mer, ger ensinnestillstånd där ingenting är omöjligt. I det ögonblick man får in i"Expert" state of mind ett stort antal saker blir omöjlig.
		-- From Henry Ford Sr., "My Life and Work"

%
Ingenting är klar förrän pappersarbetet är avklarat.
		-- From Henry Ford Sr., "My Life and Work"

%
Ingenting är omöjligt för den som inte har att göra det själv.
		-- A. H. Weiler

%
Ingenting är mer beundransvärd än mod som miljonärertolerera nackdelarna med sin rikedom.
		-- Nero Wolfe

%
Ingenting gör en person mer produktiva än i sista minuten.
		-- Nero Wolfe

%
Ingenting motiverar en man mer än att se sin chef sätta på ett ärligt dagsverke.
		-- Nero Wolfe

%
Ingenting avtar som framgång.
		-- Walter Winchell

%
Framgång föder överskott.
		-- Oscar Wilde

%
Framgång föder framgång.
		-- Alexandre Dumas

%
Framgång föder utseendet på framgång.
		-- Christopher Lascl

%
Ingenting kommer att skingra entusiasm som en liten inträdesavgift.
		-- Kim Hubbard

%
Ingenting kommer någonsin försökt om alla eventuella invändningar måste vara förstbetagen.
		-- Dr. Johnson

%
Nu kanske du frågar, "Hur kan jag få en av dessa komplett hem verktygsätter för under $ 4? "En utmärkt fråga.Gå till en av de riktigt billiga lågprisbutiker där de säljerplast möbler i färger synliga från planeten Neptunus och där dehar en del mat som specialiserat sig på pappkartonger fulla av Raisinets ochmältat mjölk bollar som tillverkats under Nixon administrationen. I enderahårdvaran eller husgeråd avdelning, hittar du ett objekt som importerats från endunkla Oriental land och beskrivs som "Nio verktyg i ett", bestående avlite handtag med utbytbara ändar representerar outgrundlig Orientalföreställningar om verktyg som amerikaner kan använda i hemmet. Köp det.Detta är den typ av verktyg som proffsen använder. Inte bara är detbillig, men det har också en stor säkerhetsfunktion som inte finns iså kallade kvalitetsverktyg set: Handtaget kommer faktiskt bryta rätt off omdu råkar slå dig själv eller något annat, eller utsätta det för direktsolljus.
		-- Dave Barry, "The Taming of the Screw"

%
Av alla möjliga utskotts reaktioner på en viss punkt på dagordningen, denreaktion som kommer att inträffa är en som kommer att frigöra den störstamängd varm luft.
		-- Thomas L. Martin

%
Naturligtvis finns det ingen anledning till det, det är bara vår politik.
		-- Thomas L. Martin

%
När den träffar fläkten, är det enda rationella val för att sopa upp, förpacka den,och sälja den som gödsel.
		-- Thomas L. Martin

%
En vacker dag, gick busschauffören att bussgarage, började sin buss,och körde iväg längs vägen. Inga problem för de första stopp - ett parmänniskor fick på, några fick, och det gick i allmänhet väl. Vid nästastopp, men en stor hulk av en kille fick på. Sex fot åtta, byggd som enbrottare, armarna hängande ner till marken. Han blängde på föraren och sade,"Big John inte betala!" och satte sig längst bak.Nämnde jag att föraren var fem fot tre, tunn, och i principödmjuk? Tja, var han. Naturligtvis gjorde han inte argumentera med Big John, men han var integlad över det. Tja, nästa dag samma sak hände - Big John fick påigen, gjorde en show att vägra att betala, och satte sig ner. Och nästa dag, ochett efter det, och så vidare. Detta riven på busschauffören, som börjadeförlora sömn över hur Big John att dra nytta av honom. slutligen hankunde stå det längre. Han undertecknade upp för bodybuilding kurser, karate, judo,och allt det bra grejer. I slutet av sommaren, hade han blivit ganska stark;vad mer, kände han riktigt bra om sig själv.Så på nästa måndag, när Big John fick återigen på bussenoch sade "Big John inte betala !," chauffören stod upp, stirrade tillbaka påpassagerare, och skrek: "Och varför inte?"Med en förvånad blick på hans ansikte, svarade Big John "Big John har enbusskort."
		-- Thomas L. Martin

%
En bra färg är värd tusen återupptas.
		-- Thomas L. Martin

%
En mans hjärna plus en annan kommer att producera en hälften så många idéer som enman skulle ha producerats enbart. Dessa två plus två mer kommer att producera halvigen så många idéer. Dessa fyra plus fyra mer börjar att representera enkreativt möte, och förhållandet ändras till en fjärdedel så många ...
		-- Anthony Chevins

%
En av dina äldsta författare, historiker vid namn Herodotos, berättar om entjuv som skulle ha verkställts. När han fördes bort han gjorde ett fynd medkungen: på ett år skulle han lära kungens favorit häst att sjungapsalmer. De andra fångarna såg tjuven sång till häst ochskrattade. "Du kommer inte att lyckas," de berättade honom. "Ingen kan."Som tjuven svarade: "Jag har ett år, och vem vet vad som kanske på den tiden. Kungen kan dö. Hästen skulle dö. Jag skulle dö.Och kanske hästen lär sig att sjunga.
		-- "The Mote in God's Eye", Niven and Pournelle

%
En möjlig orsak till att saker och ting inte går enligt planär att det aldrig fanns en plan i första hand.
		-- "The Mote in God's Eye", Niven and Pournelle

%
En lovande koncept som jag kom upp med genast var att man kundetillverkar personliga krockkuddar, sedan få en lag som antogs som kräver att de ärinstallerad på congressmen för att hålla dem från att ta resor. Låt oss säga att dinkongressledamot försökte att resa till Paris för att göra en undersöknings studie om hurden franska regeringen hanterar sjukdomar som överförs av sorbet. Just när hankom till planet, hans obligatoriska krockkudde, fastspänd runt midjan, skulleblåsa - FWWAAAAAAPPPP - vilket gör honom alltför stor för att passa genomplan dörr. Det kan också vara monterat för att blåsa upp närhelst congressmanföreslagit en lag. ( "Herr talman, folk frågar mig, varför skulle oktober varabetecknas som Cuticle besiktningsmånaden? Och jag svarar att FWWAAAAAAPPPP. ")Detta skulle spara miljontals dollar, så jag har inga tvivel om att den offentligaskulle våldsamt stödja en lag som kräver krockkuddar på kongressledamöter. Problemetär att din potentiella marknad är mycket liten: det finns bara omkring 500medlemmar av kongressen, och en del av dem, till exempel representanthusets talman "Tip" O'Neil,är redan alltför stor för att passa på normal flygplan.
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Ett sätt att göra din gamla bil köra bättre är att leta upp priset på en ny modell.
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Endast genom hårt arbete och uthållighet kan man verkligen lida.
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Möjligheter brukar förklädd till hårt arbete, så de flesta människor intekänna igen dem.
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Optimismen är innehållet i små män i höga platser.
		-- F. Scott Fitzgerald, "The Crack Up"

%
Eller du eller jag måste ge upp sitt liv till Ahrimanes. Jag skulle hellre det var du.Jag skulle inte tveka att offra mitt eget liv för att skona er, menvi tar lager nästa vecka, och det skulle inte vara rättvist mot företaget.
		-- J. Wellington Wells

%
Vår verksamhet i livet är inte att lyckas utan att fortsätta att misslyckas uppsluppen.
		-- Robert Louis Stevenson

%
Vårt land har massor av bra fem-cents cigarrer, men problemet ärde tar femton cent för dem.
		-- Robert Louis Stevenson

%
Vår policy är, när du är osäker, gör det rätta.
		-- Roy L. Ash, ex-president, Litton Industries

%
Övertrasserat? Men jag har fortfarande kontroller kvar!
		-- Roy L. Ash, ex-president, Litton Industries

%
Owe ingen något ...
		-- Romans 13:8

%
Människor är alltid tillgängliga för arbete i förfluten tid.
		-- Romans 13:8

%
Folk verkar tro att filten frasen, "Jag arbetar bara här," frikännerdem helt från någon moralisk skyldighet när det gäller allmänheten - men dettavar just Eichmanns ursäkt för sitt jobb i koncentrationslägren.
		-- Romans 13:8

%
Folk kommer att köpa något som är en till en kund.
		-- Romans 13:8

%
Vänligen hålla fingrarna borta sekreterarens reproducerande utrustning.
		-- Romans 13:8

%
Försök att begränsa mängden "detta rum inte har några bazingas"tills du blir tillsagd att dessa rum är "stansas ut." Gång utstansade,Vi har rätt att klaga illdåd, saknade bazingas, och sådant.
		-- N. Meyrowitz

%
VVS är en av de lättare av gör-det-själv-verksamhet,kräver endast några enkla verktyg och en vilja att hålla armen i enigensatt toalett. I själva verket kan du lösa många hem VVS problem, såsomirriterande kran droppa, bara genom att vrida upp radion. Men innan vi fåri specifika tekniker, låt oss titta på hur VVS fungerar.En VVS-system är mycket lik din elektriska system, med undantagatt istället för elektricitet, den har vatten, och i stället för trådar, har denrör, och i stället för radio och våffeljärn, har det kranar och toaletter.Så sanningen är att dina avlopp är ingenting alls som dinelsystem, vilket är bra, eftersom el kan döda dig.
		-- Dave Barry, "The Taming of the Screw"

%
Porsche: finns helt enkelt ingen ersättning.
		-- Risky Business

%
Ägodelar öka för att fylla det tillgängliga utrymmet för att lagra.
		-- Ryan

%
Praktiska människor skulle vara mer praktiskt om de skulle ta en litenmer tid för att drömma.
		-- J. P. McEvoy

%
Lova henne något, men ge henne Exxon blyfri.
		-- J. P. McEvoy

%
Lovande kostar ingenting, det är att leverera som dödar dig.
		-- J. P. McEvoy

%
Punktlighet är sin egen belöning, om man bor vid klockan i stället för svärdet.
		-- J. P. McEvoy

%
Sätt inte ditt förtroende i pengar, men placerar dina pengar i förtroende.
		-- J. P. McEvoy

%
Sätt din bästa fot framåt. Eller bara ringa in och säga att du är sjuk.
		-- J. P. McEvoy

%
Sätt din näsa till slipstenen!
		-- Amalgamated Plastic Surgeons and Toolmakers, Ltd.

%
Kvantitet är ingen ersättning för kvalitet, men dess enda vi har.
		-- Amalgamated Plastic Surgeons and Toolmakers, Ltd.

%
Real rikedom kan bara öka.
		-- R. Buckminster Fuller

%
Ta emot en miljon dollar skattefritt får dig att må bättre änvara pank och har ont i magen.
		-- Dolph Sharp, "I'm O.K., You're Not So Hot"

%
Nya investeringar kommer att ge en liten vinst.
		-- Dolph Sharp, "I'm O.K., You're Not So Hot"

%
Nyare forskning har tenderat att visa att den avskyvärda No-Manersätts av de dryga Procrastinator.
		-- C. N. Parkinson

%
Oavsett om ett uppdrag expanderar eller kontrakt, administrativoverhead fortsätter att växa i jämn takt.
		-- C. N. Parkinson

%
Kom ihåg - endast 10% av vad som helst kan vara i topp 10%.
		-- C. N. Parkinson

%
Kom ihåg att säga hej till din bank teller.
		-- C. N. Parkinson

%
Kom ihåg att även om du vinner rat race - du fortfarande en råtta.
		-- C. N. Parkinson

%
Pension innebär att när någon säger "Ha en bra dag", dufaktiskt har en chans på den.
		-- C. N. Parkinson

%
Riches omfattar en mängd ve.
		-- Menander

%
Regel # 7: Tystnad är inte samtycke.I motsats till vad du kanske har hört, är tystnad av de närvarandeinte nödvändigtvis samtycker, även den motvilliga sorten. De kan helt enkeltsitta i bedövas tystnad och räkna sätt att sabotera planen efterde återfår sin fattning.
		-- Menander

%
Spara lite pengar varje månad och i slutet av året kommer du attförvånad över hur lite du har.
		-- Ernest Haskins

%
Sears har allt.
		-- Ernest Haskins

%
Serverar kaffe på flygplan orsakar turbulens.
		-- Ernest Haskins

%
"Sju år och sex månader!" Humpty Dumpty upprepas tänk."En obekväm slags ålder. Nu om du hade bett mitt råd, jag skulle hasade "Lämna ut på sju" -. men det är för sent nu ""Jag ber aldrig råd om att växa," Alice sa indignerat."För stolt?" den andra frågade.Alice kände ännu mer upprörd över detta förslag. "Jag menar,"Hon sade, "att man inte kan hjälpa allt äldre.""Man kan inte, kanske", sa Humpty Dumpty; "Men två kan. Medordentlig hjälp, kanske du slutade vid sju. "
		-- Lewis Carroll, "Through the Looking-Glass"

%
För flera år sedan hade några smarta affärsmän en idé: Varför inte bygga en storbutik där en gör-det-självare kan få allt han behövde till rimligapriser? Då bestämde de sig, nah, fan med det, låt oss bygga ett hemcentrum. Och snart hem centra växer upp som crabgrass allaöver hela USA.
		-- Dave Barry, "The Taming of the Screw"

%
Visa mig en människa som är en god förlorare och jag ska visa dig en man som spelargolf med sin chef.
		-- Dave Barry, "The Taming of the Screw"

%
Så du tror att pengar är roten till allt ont. Har du någonsin frågat vadär roten till pengarna?
		-- Ayn Rand

%
Så ... har du någonsin undrar, gör garbagemen ta duschar innan de går till jobbet?
		-- Ayn Rand

%
Vissa människor rista karriärer, andra mejsel dem.
		-- Ayn Rand

%
Vissa människor har en stor ambition: att bygga någotsom kommer att pågå åtminstone tills de är färdiga med att bygga det.
		-- Ayn Rand

%
Vissa människor hantera genom boken, trots att de inte vet vem skrevbok eller ens vilken bok.
		-- Ayn Rand

%
Vissa människor bara öppna upp för att berätta att de är stängda.
		-- Ayn Rand

%
Vissa människor ber för mer än vad de är villiga att arbeta för.
		-- Ayn Rand

%
Vissa människor säger en frontmotor bil hanterar bäst. Vissa människor säger enbak-motor bil hanterar bäst. Jag säger en hyrd bil hanterar bäst.
		-- P. J. O'Rourke

%
Någon borde korsa kulspetspennor med galgar så attpennor kommer att öka i stället för att försvinna.
		-- P. J. O'Rourke

%
Någon gång i framtiden någon har fått för att avgöra om skrivmaskinen är maskinen,eller den person som driver det.
		-- P. J. O'Rourke

%
Someday utskrifterna kommer.
		-- Kodak

%
Någon är unenthusiastic om ditt arbete.
		-- Kodak

%
Suburbia är där utvecklaren bulldozes ut träden, sedan namngatorna efter dem.
		-- Bill Vaughn

%
Framgång är något jag kommer att klä sig för när jag kommer dit, och inte förrän.
		-- Bill Vaughn

%
Föreslår du bara sitta där och vänta tills livet blir lättare.
		-- Bill Vaughn

%
Stötta din lokala kyrka eller synagoga. Bedja vid Bank of America.
		-- Bill Vaughn

%
Överraskning förfaller idag. Även hyran.
		-- Bill Vaughn

%
Överraska din chef. Få tid till jobbet.
		-- Bill Vaughn

%
Ta hand om lyx och förnödenheter kommer att ta hand om sig själva.
		-- Lazarus Long

%
Ta allt i steg. Trampa alla som kommer i din väg.
		-- Lazarus Long

%
Ta folks vid Coca-Cola. Under många år var de innehållatt luta sig tillbaka och göra samma gamla kolsyrad dryck. Det var en bradryck, ingen tvekan om det, generationer av människor hade vuxit uppdricka det och göra experiment i sexan där du sätter enspika i ett glas av koks och efter ett par dagar spik löser uppoch läraren säger: "Tänk vad det gör att tänderna!" Så Coca-Colavar stabilt förankrade på marknaden, och ledningen såg inget behov av attförbättra ...
		-- Dave Barry, "In Search of Excellence"

%
Ta dig tid att reflektera över alla de saker du har, inte som ett resultat av dinförtjänst eller hårt arbete eller på grund av Gud eller slumpen eller insatser för andra människorhar gett dem till dig.
		-- Dave Barry, "In Search of Excellence"

%
Ta ditt arbete på allvar men aldrig ta sig själv på allvar; och inteta vad som händer antingen själv eller ditt arbete på allvar.
		-- Booth Tarkington

%
Talang gör vad den kan.Genius gör vad den måste.Du gör vad du får betalt för att göra.
		-- Booth Tarkington

%
Telefonkataloger är som ordböcker - om du vet svaret innandu slå upp det, kan du så småningom bekräftar vad du trodde du visstemen var inte säker. Men om du söker efter något som du interedan vet, fingrarna kunde gå själva till döds.
		-- Erma Bombeck

%
Term, helgdagar, term, helgdagar, tills vi lämnar skolan, och sedan arbeta, arbete,arbeta tills vi dör.
		-- C. S. Lewis

%
Sånt är livet.Vad är livet?En tidning.	Hur mycket kostar det?Två-fifty.Jag har bara en dollar.Sånt är livet.
		-- C. S. Lewis

%
Den [Ford Foundation] är en stor mängd pengar helt omgiven avmänniskor som vill ha lite.
		-- Dwight MacDonald

%
Det så kallade ensamvarg "kan respekteras, men han är alltid förbittrade av hans kollegor,för han verkar vara passerar en kritisk bedömning av dem, när han kan varahelt enkelt göra en begränsande uttalande om sig själv.
		-- Sidney Harris

%
Frånvarande som är alltid fel.
		-- Sidney Harris

%
Svaret på frågan om livet, universum och allt är ...Fyra dagars arbetsvecka,Två skikt toalettpapper!
		-- Sidney Harris

%
Svaret på den ultimata fråga om liv, universum och allt varsläpps med tillstånd av Amalgamated unionen filosofer,Vise, armatur, och andra professionella tänkande personer.
		-- Sidney Harris

%
Den genomsnittliga individens ställning i någon hierarki är mycket som att drahundspann - det finns ingen verklig miljöombyte med undantag för ledarhund.
		-- Sidney Harris

%
Den bästa utrustningen för ditt arbete är naturligtvis den dyraste.Dock är din granne alltid slösa pengar som borde vara dingenom att bedöma saker vid deras pris.
		-- Sidney Harris

%
Den bästa verkställande är en som har förstånd nog att plocka goda människor att göravad han vill ha gjort, och självbehärskning tillräckligt för att hålla från inblandning meddem medan de gör det.
		-- Theodore Roosevelt

%
De bästa som planer på möss och män hålls upp i den juridiska avdelningen.
		-- Theodore Roosevelt

%
De bästa sakerna i livet är mot en avgift.
		-- Theodore Roosevelt

%
De bästa sakerna i livet att börja säljas förr eller senare.
		-- Theodore Roosevelt

%
Det bästa sättet att undvika ansvar är att säga, "Jag har ansvar."
		-- Theodore Roosevelt

%
Bibeln på bokstäverna i referens:Börjar vi om igen för att producera våra referenser? Dovi, som vissa människor behöver introduktionsbrev till dig, eller från dig?Nej, du är alla brev vi behöver ett brev skrivet på ditt hjärta; någraman kan se det för vad det är och läsa det för sig själv.
		-- 2 Corinthians 3:1-2, New English translation

%
Det största misstaget du kan göra är att tro att du arbetar förnågon annan.
		-- 2 Corinthians 3:1-2, New English translation

%
Chefen återvänt från lunch på gott humör och kallade hela personalenför att lyssna på ett par skämt han hade plockat upp. Alla utom en flickaskrattade uproariously. "Vad är problemet?" muttrade chefen. "Har du intefick en känsla för humor? ""Jag behöver inte skratta", sade hon. "Jag lämnar fredag ​​ändå.
		-- 2 Corinthians 3:1-2, New English translation

%
Hjärnan är en underbar organ; det börjar arbeta så fort du får upppå morgonen, och inte sluta förrän du kommer till jobbet.
		-- 2 Corinthians 3:1-2, New English translation

%
Den närmaste till perfektion en person någonsin kommer är när han fyller ut ett jobbansökningsblankett.
		-- Stanley J. Randall

%
Förvirringen av en anställd mäts genom längden på sina minnesanteckningar.
		-- New York Times, Jan. 20, 1981

%
Kostnaden för fjädrar har ökat, även ner är upp!
		-- New York Times, Jan. 20, 1981

%
Levnadskostnaderna har inte påverkat dess popularitet.
		-- New York Times, Jan. 20, 1981

%
Levnadskostnaderna går upp, och chansen att leva går ner.
		-- New York Times, Jan. 20, 1981

%
Beslutet behöver inte vara logiskt; Det var enhälligt.
		-- New York Times, Jan. 20, 1981

%
Graden av teknisk förtroende är omvänt proportionell mot denledningsnivå.
		-- New York Times, Jan. 20, 1981

%
Den avgående division general manager träffade en sista gång med sin ungaefterträdare och gav honom tre kuvert. "Min företrädare gjorde detta för mig,och jag kommer att passera traditionen vidare till dig ", sade han." Vid första teckenproblem, öppna det första kuvertet. Eventuella ytterligare svårigheter, öppnaandra höljet. Sedan, om problemen fortsätter, öppna den tredje kuvertet.Lycka till. "Den nya chefen återvände till sitt kontor och kastade kuverteni en låda.Sex månader senare, kostnader skjutit i höjden och resultatet rasade. Skakad, denung man öppnade första kuvertet, som sagt, "skylla allt på mig."Nästa dag, höll han en presskonferens och gjorde just detta. Dekris passerade.Sex månader senare, minskade försäljningen tvärt. belägradechef öppnade andra kuvertet. Det sade, "Omorganisera."Han höll en annan presskonferens och meddelade att uppdelningenskulle omstruktureras. Krisen passerat.Ett år senare, allt gick fel på en gång och chefen varskulden för allt. Den härjade verkställande stängde sitt kontor dörr, sjönki sin stol, och öppnade tredje kuvertet."Förbered tre kuverten ..." det sagt.
		-- New York Times, Jan. 20, 1981

%
Skillnaden mellan en karriär och ett jobb är cirka 20 timmar per vecka.
		-- New York Times, Jan. 20, 1981

%
Den svåra vi gör idag; det omöjliga tar lite längre tid.
		-- New York Times, Jan. 20, 1981

%
Early bird som fångar masken fungerar för någon som kommer i slutet avoch äger masken gården.
		-- Travis McGee

%
Det enklaste sättet att räkna levnadskostnaderna är att ta dina inkomster ochlägga tio procent.
		-- Travis McGee

%
I slutet av arbetskraft är att få fritid.
		-- Travis McGee

%
Felet ungdomar är att tro att intelligens är ett substitut förerfarenhet, medan felet ålder är att tro erfarenhet är ett substitutför intelligens.
		-- Lyman Bryson

%
Ju snabbare jag går, den behinder jag får.
		-- Lewis Carroll

%
Den finaste vältalighet är det som får saker och ting gjorda.
		-- Lewis Carroll

%
Den första 90% av ett projekt tar 90% av tiden, tar den sista 10% avövriga 90% av tiden.
		-- Lewis Carroll

%
Den första myten om ledningen är att det existerar. Den andra myten omförvaltning är att framgång är lika med skicklighet.
		-- Robert Heller

%
Den första rotarian var den förste att kalla Johannes Döparen "Jack".
		-- H. L. Mencken

%
Den första regeln av intelligent mixtrande är att spara alla delar.
		-- Paul Erlich

%
Den vattentoalett är grunden för den västerländska civilisationen.
		-- Alan Coult

%
Gent som vaknar upp och befinner sig en framgång har inte sovit.
		-- Alan Coult

%
Den största produktivkraft är människans själviskhet.
		-- Robert Heinlein

%
Den svåraste delen av klättra på stegen till framgång är att få igenompubliken längst ner.
		-- Robert Heinlein

%
Hieroglyferna är alla oläslig utom för en notering på baksidan,som lyder "Äkta äkta egyptisk papyrus. Garanterad att varaminst 5000 år gammal. "
		-- Robert Heinlein

%
Tanken var att konsumenterna skulle ta med brutna elektroniskaenheter, t.ex. TV-apparater och videobandspelare, till centra förstöring,där utbildad personal skulle döda dem (enheter) med släggor.Med sina enheter därmed permanent förstörd, skulle konsumenterna sedan vara friatt gå ut och köpa nya enheter, snarare än att slarva bort år avderas liv försöker ha de gamla repareras så kallade "fabrikservicecenter ", som i själva verket består av två män som heter Lester peta påinsidan av trasiga elektroniska apparater med billiga cigarrer och gå,"Lookit alla dem trådar i det!"
		-- Dave Barry, "'Mister Mediocre' Restaurants"

%
Den idealiska rösten för radio kan definieras som visar inget ämne, inget sex,ingen ägare och ett budskap om vikten för varje hemmafru.
		-- Harry V. Wade

%
Tomgångs man inte vet vad det är att njuta av resten.
		-- Harry V. Wade

%
Den individuella val av kvarstad av en hamburgare kan vara en viktigpekar till konsumenten i denna dag när individualism är en alltviktiga för människor.
		-- Donald N. Smith, president of Burger King

%
Intelligens varje diskussion minskar med kvadraten påantal deltagare.
		-- Adam Walinsky

%
IQ gruppen är den lägsta IQ av en medlem av gruppen delasmed antalet personer i gruppen.
		-- Adam Walinsky

%
Kungen och hans rådgivare har utsikt över slagfältet:King: "Hur går stridsplan?"Handledare: "Se dessa små svarta prickar som kör till höger?"K: "Ja."A: "De är deras killar och alla dessa små röda prickar igång.till vänster är våra killar. Sedan när de kolliderar vi vänta tillsdammet försvinner. "K: "Och"A: "Om det finns fler röda fläckar kvar än svarta fläckar, vinner vi."K: "Men hur är det ^ # !! $% stridsplan?"A: "Hittills verkar det att gå enligt fläckar."
		-- Adam Walinsky

%
Den sista personen som slutade eller fick sparken kommer att hållas ansvariga förallt som går fel - tills nästa person avslutas eller bränns.
		-- Adam Walinsky

%
Ju längre titeln, den mindre viktig jobbet.
		-- Adam Walinsky

%
Den stora skillnaden mellan obligationer och obligationshandlare är att obligationerna kommersmåningom mogna.
		-- Adam Walinsky

%
Medlet-och-slutar moralister, eller icke-doers, alltid hamnar på deras ändarutan något sätt.
		-- Saul Alinsky

%
De ödmjuka vill inte ha den.
		-- Saul Alinsky

%
De ödmjuka skall ärva jorden - de är för svaga för att vägra.
		-- Saul Alinsky

%
De ödmjuka skall ärva jorden, men * inte * sina rättigheter mineral.
		-- J. P. Getty

%
De ödmjuka skall ärva jorden. (Men de kommer att kämpa för det.)
		-- J. P. Getty

%
De ödmjuka skall ärva jorden; men då det inte kommer att varanågot kvar värt ärva.
		-- J. P. Getty

%
Desto mer hjärtlig köparens sekreterare, desto större är oddsen att denkonkurrens har redan ordern.
		-- J. P. Getty

%
Ju mer skit du stå ut med, desto mer skit du ska få.
		-- J. P. Getty

%
Ju mer jag vill få något gjort, ju mindre jag kallar det att fungera.
		-- Richard Bach, "Illusions"

%
Ju mer pretentiös ett företags namn, desto mindre organisationen. (FörExempelvis Murphy Center för kodifiering av mänsklig och organisatorisk lag,kontrast till IBM, GM, AT & T ...)
		-- Richard Bach, "Illusions"

%
Den mest härlig dag efter den på vilken du köper en stuga ilandet är en som du sälja den.
		-- J. Brecheux

%
Det svåraste i världen är att veta hur man gör en sak och atttitta på någon annan gör det fel, utan att kommentera.
		-- T. H. White

%
En dag du vill sälja din själ för något, själar är ett överflöd.
		-- T. H. White

%
Det enda problemet med att vara en man av fritid är att man aldrig kan slutaoch ta en paus.
		-- T. H. White

%
De enda främjande regler jag kan komma på är att en känsla av skam är attundvikas till varje pris och det finns aldrig någon anledning till en hustler tillvara mindre listig än mer dygdiga män. Oh ja ... när du trordu har något riktigt bra, lägga till tio procent mer.
		-- Bill Veeck

%
Den enda riktigt bra ställe att köpa virke är en butik där virket harredan skurits och fästs samman i form av möbler, färdiga,och sätta in lådor.
		-- Dave Barry, "The Taming of the Screw"

%
Opossumen är en mycket sofistikerad djur. Det behöver inte ens få upptills 5 eller 6:00.
		-- Dave Barry, "The Taming of the Screw"

%
Den optimala kommitté har inga medlemmar.
		-- Norman Augustine

%
Överflöd av front office dörren varierar omvänt med den fundamentalasolvens företaget.
		-- Norman Augustine

%
Den andra raden flyttas snabbare.
		-- Norman Augustine

%
Den person som kan le när något går fel har tänkt pånågon att skylla det på.
		-- Norman Augustine

%
Den person som gör inga misstag brukar inte göra någonting.
		-- Norman Augustine

%
Den person som tar dig till lunch har inte för avsikt att betala.
		-- Norman Augustine

%
Innehav av en bok blir ett substitut för att läsa det.
		-- Anthony Burgess

%
Priset man betalar för att uppnå något yrke, eller ringa, är en intimkunskap om sitt fula sida.
		-- James Baldwin

%
Den primära orsaken till fel i elektriska apparater är ett utgångetgaranti. Ofta kan du få en apparat igång igen bara genom att ändragarantiutgångsdatum med en 15/64 tum filtmarkör.
		-- Dave Barry, "The Taming of the Screw"

%
Det problem som vi trodde var ett problem var verkligen ett problem, meninte problemet vi trodde var problemet.
		-- Mike Smith

%
Anledningen till oron dödar fler människor än arbete är att fler människororoa än arbete.
		-- Mike Smith

%
Belöningen för att arbeta hårt är mer hårt arbete.
		-- Mike Smith

%
Belöningen för en sak bra gjort är att ha gjort det.
		-- Emerson

%
De rika blir rika och fattiga blir fattigare.De rika får mer, de som inte har dö.
		-- Emerson

%
Rättigheter och intressen arbetande mannen kommer att skyddas och vårdasför att inte våra arbets agitatorer, men de kristna män som Gud i sinoändliga visdom har gett kontroll av egendom intressen i landet, ochpå framgångsrik förvaltning som så mycket som återstår.
		-- George F. Baer, railroad industrialist

%
Vägen till undergång är alltid i gott skick, och de resenärerna betalabekostnad av den.
		-- Josh Billings

%
Lönen för verkställande av stort företag är inte en marknadPriset för prestation. Det är ofta i form av en varm personliggest av individen själv.
		-- John Kenneth Galbraith, "Annals of an Abiding Liberal"

%
Hemligheten bakom framgången är uppriktighet. När du kan falska att du hardet gjorde.
		-- Jean Giraudoux

%
De sju dödssynderna ... Mat, kläder, bränning, hyra, skatter, respektabilitetoch barn. Ingenting kan lyfta dessa sju milstolpar från mannens hals menpengar; och ande kan inte sväva förrän milstolparna lyfts.
		-- George Bernard Shaw

%
Det kortaste avståndet mellan två punkter är under uppbyggnad.
		-- Noelie Alito

%
Ju tidigare du halkar efter, desto mer tid du har att komma ikapp.
		-- Noelie Alito

%
Ju tidigare du gör din första 5000 misstag, desto snabbare kommer du attkunna rätta till dem.
		-- Nicolaides

%
Stjärnan i rikedom skiner på dig.
		-- Nicolaides

%
Den överlägsna mannen förstår vad som är rätt; sämre man förstårvad kommer att sälja.
		-- Confucius

%
Termen "eld" tar upp visioner av våld och förödelse och fula scenenskytte medarbetare som gör misstag. Vi kommer nu att hänvisa till denna processsom "ta bort" en anställd (mycket som en fil tas bort från en disk). Deanställd är helt enkelt det ett ögonblick, och borta nästa. All den fruktansvärdavredesutbrott, gråt, och hot elimineras.
		-- Kenny's Korner

%
Tiden på någon punkt på dagordningen [av ett finansutskott] kommer att varai omvänd proportion till den berörda summan.
		-- C. N. Parkinson

%
Problemet med en hel del självgjorda män är att de dyrkar sin skapare.
		-- C. N. Parkinson

%
Problemet med att vara fattig är att det tar upp all din tid.
		-- C. N. Parkinson

%
Problemet med att vara punktliga är att ingen är där för att uppskatta det.
		-- Franklin P. Jones

%
Problemet med att vara punktliga är att folk tror att du har inget merviktigt att göra.
		-- Franklin P. Jones

%
Problemet med att göra något rätt första gången är att ingenuppskattar hur svårt det var.
		-- Franklin P. Jones

%
Problemet med pengar är det kostar för mycket!
		-- Franklin P. Jones

%
Problemet med möjlighet är att det alltid kommer förklädd till hårt arbete.
		-- Herbert V. Prochnow

%
Problemet med ekorrhjul är att även om du vinner, du är fortfarande en råtta.
		-- Lily Tomlin

%
De två mest vackra ord i det engelska språket är "Check Länkade."
		-- Dorothy Parker

%
Användningen av pengar är all fördel finns att ha pengar.
		-- B. Franklin

%
Syndens lön är hög men du får dina pengar värde.
		-- B. Franklin

%
Syndens lön är orapporterat.
		-- B. Franklin

%
Sättet att göra en liten förmögenhet på råvarumarknaden är att börjamed en stor förmögenhet.
		-- B. Franklin

%
Den värsta biluthyrningNär David Schwartz lämnade universitetet i 1972, satte han upp Rent-A-Wrecksom ett skämt. Att vara en naturlig upptågsmakare, fick han en flotta av beat-upsjaskigt, wreckages väntar på skrothögen i Kalifornien.Han satte på ett lock och såg fram emot att titta på människors ansikten som hanförde dem runt valet av bumperless, bucklade junkmobiles.Till sin varaktig förvåning var en omättlig efterfrågan på dem ochHan har nu 26 blomstrande filialer över hela Amerika. "Folk gillar körningrunda i värsta bilar tillgängliga ", sade han. Naturligtvis de gör."Om föraren skadar sidan av en bil och är ärliga nog atterkänna det, säger jag honom: 'Glöm det. Om de tar en bil tillbaka sent viförbise det. Om de har haft en krasch och det innebär inte ett annat fordonvi kan bortse från det också. ""Var är askkoppen?" frågade en Los Angeles fru, som hon fasti de rippade interiören. "Älskling", sa hennes man, "hela bilen äraska fack. "
		-- Stephen Pile, "The Book of Heroic Failures"

%
Deras idé om ett erbjudande du inte kan vägra är ett erbjudande ... och du är bästinte vägra.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Dem som har, blir.
		-- Stephen Pile, "The Book of Heroic Failures"

%
Då sade en man: Prata med oss ​​av förväntningar.Han sade då: Om en man inte se eller höra vattenJordanien, då han ska inte smaka granatäpple eller ply sina varor i enöppen marknad.Om en människa skulle inte arbete i salt och bergtäkter sedan hanbör inte acceptera av jorden det som han vägrar att ge avhan själv.En sådan man skulle förvänta sig ett päron av en persika träd.En sådan man skulle förvänta sig en sten för att lägga ett ägg.En sådan man skulle förvänta sig Sears att montera en gräsklippare.
		-- Kehlog Albran, "The Profit"

%
Sedan fanns det Scoutmasteren som fick en fantastisk affär på detta fallTates varumärke kompasser för hans troup; endast $ 1.25 varje! Enda problemet var,när de fick dem ut i skogen, de kompasser var alla fastnat pekartill "W" på ratten.Moralisk:Den som har en Tates är förlorad!
		-- Kehlog Albran, "The Profit"

%
Det finns många av oss i denna gamla världen till oss som menar att saker går sönderom även för oss alla. Jag har observerat, till exempel, att vi alla fårungefär samma mängd av is. De rika blir det på sommaren och de fattigafå det på vintern.
		-- Bat Masterson

%
Det finns värre saker i livet än döden. Har du någonsin tillbringat en kvällmed en försäkring försäljare?
		-- Woody Allen

%
Det har varit lite nöd sälja på börsen.
		-- Thomas W. Lamont, October 29, 1929 (Black Tuesday)

%
Det finns en hel del högtidlig cant om gemensamma intressen kapitaloch arbetskraft. Som det står, är deras enda gemensamma intresse att skärvarandras hals.
		-- Brooks Atkinson, "Once Around the Sun"

%
Det finns knappast en sak i världen att någon man inte kan göra en litensämre och sälja lite billigare.
		-- Brooks Atkinson, "Once Around the Sun"

%
Det finns aldrig tid att göra det rätt, men alltid tid att göra det.
		-- Brooks Atkinson, "Once Around the Sun"

%
"Det finns ingen jultomten. Det är bara en marknadsföring knep för att göra låg inkomstföräldrars liv ett elände. ""... Jag vill att du ska föreställa lita ett barns ansikte, strimmig med tårarpå grund av vad du just sa. ""Jag vill att du ska föreställa ansiktet på sin mor, eftersom en veckas Dole kommer intebetala för en Master of the Universe Jagare! "
		-- Filthy Rich and Catflap

%
Det finns ingen tid som den nuvarande för att skjuta upp vad du borde göra.
		-- Filthy Rich and Catflap

%
Det finns inget så lätt, men att det blir svårt när du gör detmotvilligt.
		-- Publius Terentius Afer (Terence)

%
Det är ett sätt att ta reda på om en man är ärlig - fråga honom. Om han säger"Ja" du vet att han är krokig.
		-- Groucho Marx

%
Det finns mycket lite framtid att vara rätt när din chef är fel.
		-- Groucho Marx

%
Det måste finnas mer i livet än att ha allt.
		-- Maurice Sendak

%
Det fanns en högskolestudent försöker tjäna lite fickpengar genomgå från hus till hus erbjudande att göra udda jobb. Han förklarade detta fören man som svarade en dörr."Hur mycket kommer du ladda att måla min veranda?" frågade mannen."Fyrtio dollar.""Fine" sade mannen, och gav studenten färg och penslar.Tre timmar senare paint-stänkte lad knackade på dörren igen."Klart!", Säger han, och samlar sina pengar. "Förresten," eleven säger"Det är inte en Porsche, det är en Ferrari."
		-- Maurice Sendak

%
Det finns inget sådant som en gratis lunch.
		-- Milton Friendman

%
Det finns inget värre för din verksamhet än extra jultomtarrökning i män rum.
		-- W. Bossert

%
De är dårar som tror att rikedom eller kvinnor eller starka drycker eller ensdroger kan köpa det mesta i försök av själen i en människa. Dessa saker harbleka nöjen jämfört med det som är störst av dem alla, sitt uppdrag, somkrav från honom mer än sitt yttersta styrka, absorberar honom att, ben ochmuskel och hjärna och hopp och rädsla och drömmar - och ändå kräver mer.De är dårar som tror något annat. Inga stora ansträngningar någonsin köpt.Ingen målning, ingen musik, ingen dikt, ingen katedral i sten, ingen kyrka, ingen stat varnågonsin höjs till stånd för betalning av något slag. Ingen parthenon, ingen Thermopylaenågonsin byggts eller kämpat för lön eller ära; ingen Bukhara sparken, eller Kina markunder Mongol häl, för byte eller makt ensam. Betalningen för att göra dessasaker var själv göra av dem.Svinga sig - att använda sig själv som ett verktyg i den egna sidan - ochså att göra eller bryta det som ingen annan kan bygga eller förstöra - det ärstörsta nöje som människan känner till! Till en som har känt mejseln i handenoch befria ängeln fängslad i marmorblocket, eller en som har käntsvärd i handen och ställa hemlösa själen som en stund innan bodde i kroppenav hans dödsfiende - till dem båda kommer både smaken av den sällsynta matspridas endast för demoner eller gudar. "
		-- Gordon R. Dickson, "Soldier Ask Not"

%
Saker värt att ha är värt att fuska för.
		-- Gordon R. Dickson, "Soldier Ask Not"

%
Tänk tur. Om du faller i en damm, kontrollera dina fickor för fisk.
		-- Darrell Royal

%
Detta är ett bra tillfälle att punt arbete.
		-- Darrell Royal

%
Detta är en särskilt bra tid för dig turister som planerar att flyga, eftersomReagan-administrationen, som en del av samma politik enligt vilken detnyligen sålt Yellowstone National Park till Wayne Newton har "avreglerade"flygbranschen. Vad detta innebär för dig, konsumenten, är attflygbolagen inte längre behövs för att följa några regler alls. Dom kanvisa snuff movies. De kan ta betalt för syre. De kan hyra piloter rättav Varuautomat Refill Person School. De kan spara bränsle genomutstötning husky passagerare över vatten. De kan ramma konkurrerande plan ii luften. Dessa innovationer har lett till enorma kostnadsbesparingar somhar gått vidare till dig, konsumenten, i form av flyg medotroligt låga priser, såsom $ 29. Naturligtvis behöver vissa begränsningar,det viktigaste är att alla dessa flygningar tar dig till Newark, och du måstebetala tusentals dollar om du vill flyga tillbaka ut.
		-- Dave Barry, "Iowa -- Land of Secure Vacations"

%
Denna planet har - eller snarare hade - ett problem, som var detta: de flesta avde människor som lever på det var olycklig för ganska mycket av tiden. Mångalösningar föreslagits för detta problem, men de flesta av dessa vartill stor del sysslar med rörelser små gröna papperslappar,vilket är märkligt eftersom på det hela taget var inte de små gröna bitar avpapper som var missnöjda.
		-- Douglas Adams

%
Den här veckan bara, alla våra fiber fylla jackor markeras!
		-- Douglas Adams

%
De som hävdar de döda aldrig återvända till livet har aldrig funnitshär på avsluta tid.
		-- Douglas Adams

%
De som gör saker i en ädel anda av självuppoffring ska kunna undvikastill varje pris.
		-- N. Alexander.

%
Tid är det mest värdefulla man kan spendera.
		-- Theophrastus

%
Dags att ta lager. Gå hem med några kontorsmateriel.
		-- Theophrastus

%
För att undvika kritik, gör ingenting, säger ingenting, vara ingenting.
		-- Elbert Hubbard

%
Att vara eller inte vara, det är den nedersta raden.
		-- Elbert Hubbard

%
För att göra ingenting är att vara ingenting.
		-- Elbert Hubbard

%
Att göra två saker samtidigt är att göra heller.
		-- Publilius Syrus

%
För att komma tillbaka på fötterna, missar två bil betalningar.
		-- Publilius Syrus

%
Att få något gjort, bör en kommitté bestå av mer än trepersoner, två av dem frånvarande.
		-- Publilius Syrus

%
För att återställa en känsla av verklighet, tror jag Walt Disney skulle ha en Hardluckland.
		-- Jack Paar

%
För att spara en enda liv är bättre än att bygga en sju våningar pagod.
		-- Jack Paar

%
Att se ett behov och väntar på att bli tillfrågad, är att redan vägra.
		-- Jack Paar

%
Att upptäcka expert, välja den som förutspår jobbet tar längstoch kostar mest.
		-- Jack Paar

%
Att stanna ungdomlig, bo bra.
		-- Jack Paar

%
Till hyresvärden tillhör de dörrhandtag.
		-- Jack Paar

%
Till ditt eget själv vara sant. (Om inte det, åtminstone göra några pengar.)
		-- Jack Paar

%
För att förstå denna viktiga historia, måste man förstå hur telefonenFöretaget arbetar. Telefonen är ansluten till en lokal dator, vilket är isin tur är ansluten till en regional dator, som i sin tur är ansluten till enhögtalaren storleken av en sopbil på gräsmattan i Edna A. Bargewater avLawrence, Kan.När du talar i telefon, lyssnar din lokala dator i. Om detmisstänker att du kommer att diskutera en intim ämne, meddelar det datornovan, som lyssnar på och beslutar om att varna en ovanför,tills slutligen, om du verkligen förödmjuka dig, kanske bryta ner i tåraroch berätta för din närmaste vän om en smutsig incident från ditt förflutnainbegriper en förslappad Motell, en granne make, en hel religiös ordning, enträdgårdsslang och sex liter tapiokapudding matar top dator dinsamtal till Ednas högtalare, och hon och hennes vänner komma ut påveranda att lyssna och dricka gin och skratta sig dum.
		-- Dave Barry, "Won't It Be Just Great Owning Our Own Phones?"

%
Alltför många människor tänker på säkerhet i stället för möjligheter. De verkarmer rädd för livet än döden.
		-- James F. Byrnes

%
För mycket är inte tillräckligt.
		-- James F. Byrnes

%
För mycket av allt är precis tillräckligt.
		-- Bob Wier

%
Sanningen är gratis, men informationen kostar.
		-- Bob Wier

%
Två kan leva så billigt som en för hälften så lång.
		-- Howard Kandel

%
Veni Vidi, VISA:Jag kom, jag såg, jag gjorde lite shopping.
		-- Howard Kandel

%
Mycket få saker faktiskt få tillverkas i dessa dagar, eftersom enoändligt stora universum, som den som vi lever i, det mesta enskulle kunna tänka sig, och en hel del saker som man helst inte, växernågonstans. En skog upptäcktes nyligen i de flesta av träden växtespärr skruvmejslar som frukt. Livscykeln för den hylsmejsel ärganska intressant. När plockas det behöver en mörk dammiga låda där det kanligga ostörd i flera år. Sedan en natt plötsligt luckor, kasserar sinyttre hud som smular in damm, och framstår som en helt oidentifierbaralite metall objekt med flänsar i båda ändar och en sorts ås och ett hålför en skruv. Detta då hittas kommer kastas bort. Ingen vet vadskruvmejsel är tänkt att vinna på detta. Natur, i sin oändliga visdom,är förmodligen arbetar på det.
		-- Howard Kandel

%
Västar ska kostymer som säkerhetsbälten är bilar.
		-- Howard Kandel

%
VI:En hungrig hund jagar bäst.En hungrigare hund jagar ännu bättre.VII:Minskad affärsbasen ökar overhead.Så gör ökad affärs bas.VIII:De misslyckade fyra år i utbildningen av en kostnads ​​estimatornär femman aritmetik.IX:Akronymer och förkortningar ska användas i största möjliga utsträckningmöjligt att göra triviala idéer djupgående. Quod erat demonstrandumX:Tjurar inte vinna tjurfäktningar; människor gör.Människor inte vinner människor slagsmål; advokater gör.
		-- Norman Augustine

%
Vital papper kommer att visa sin vitalitet genom spontant flyttafrån där du lämnade dem till där du inte kan hitta dem.
		-- Norman Augustine

%
VARNING all personal:Skjutningar kommer att fortsätta tills moral förbättras.
		-- Norman Augustine

%
Avfall inte få din budget skär nästa år.
		-- Norman Augustine

%
Vi vill alla beröm, men en vandring i vår lön är den bästa sortens sätt.
		-- Norman Augustine

%
Vi lever i ett tillstånd av ambitiös fattigdom.
		-- Decimus Junius Juvenalis

%
Vi är inte en älskad organisation, men vi är en respekterad man.
		-- John Fisher

%
Vi har några helt ovedersägliga statistik för att visa exakt varfördu är så trött.Det finns inte så många människor som faktiskt arbetar som du kanske trodde.Befolkningen i det här landet är 200 miljoner. 84 miljoner är över60 år, vilket lämnar 116 miljoner för att göra jobbet. Personer under 20år totalt 75 miljoner, vilket lämnar 41 miljoner för att göra jobbet.Det finns 22 miljoner som är anställda av regeringen, som lämnar19 miljoner för att göra jobbet. Fyra miljoner är i de väpnade styrkorna, somlämnar 15 miljoner för att göra jobbet. Dra av 14.800.000, antalet i tillståndetoch stadskontor, lämnar 200.000 för att göra jobbet. Det finns 188 tusen isjukhus, mentalsjukhus, etc., så som lämnar 12000 att göra arbetet.Nu kan det intressera dig att veta att det finns 11,998 personer i fängelse,så som lämnar bara två personer för att bära lasten. Det är du och jag, ochbror, jag börjar bli trött på att göra allt själv!
		-- John Fisher

%
"Vi hävdar att själva grunden för vårt sätt att leva är vad vi kallarfri företagsamhet ", säger Cash McCall", men när en av våra medborgarevisar tillräckligt fri företagsamhet att stapla upp lite av denna vinst, vi görvårt bästa för att få honom att känna att han borde skämmas över sig själv. "
		-- Cameron Hawley

%
Vi var så dålig att vi trodde nya kläder innebar någon hade dött.
		-- Cameron Hawley

%
Vi var så dålig att vi inte kunde råd med en vakthund. Om vi ​​hörde ett ljud på natten,vi skulle skälla oss.
		-- Crazy Jimmy

%
Vi lever i en guldålder. Allt du behöver är guld.
		-- D. W. Robertson.

%
Weekend, var är du?
		-- D. W. Robertson.

%
Hur bra är en biljett till det goda livet, om du inte kan hitta ingången?
		-- D. W. Robertson.

%
Vad jag menar (och alla andra medel) med ordet kvalitet kan inte varadelas upp i ämnen och predikat. Detta beror inte på kvalitetär så mystisk men eftersom kvaliteten är så enkel, omedelbar och direkt.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad är värt att göra är värt besväret att be någon att göra.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad synd inte har begåtts i effektivitetens namn?
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad stort tryck giver, tager det finstilta bort.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad de sa:Vad de menade:"Jag rekommenderar denna kandidat med några som helst kvalifikationer."(Ja, det om sammanfattar det.)"Mängden av matematik hon vet kommer att överraska dig."(Och jag rekommenderar att du inte ger den skolan en dime ...)"Jag kan inte säga tillräckligt bra saker om honom."(Vad en skruv-up.)"Jag är glad att kunna säga att denna kandidat är en före detta kollega till mig."(Jag kan inte säga hur glad jag är att hon lämnade vårt företag.)"När den här personen lämnade vår anställa, var vi ganska hoppfull att han skulle gålångt med sina kunskaper. "(Vi hoppades att han skulle gå så långt som möjligt.)"Du kommer inte hitta många människor som henne."(I själva verket kan de flesta människor inte stå att vara omkring henne.)"Jag kan inte rekommendera honom alltför mycket."(Men, såvitt jag vet, han har aldrig begått ettbrott i min närvaro.)
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad de sa:Vad de menade:"Om du visste denna person samt jag känner honom, skulle du tänka så mycketav honom som jag gör. "(Eller så lite, att formulera det lite mer exakt.)"Hennes ingång var alltid kritisk."(Hon hade aldrig ett gott ord att säga.)"Jag har inga tvivel om hans förmåga att göra ett bra arbete."(Och det är obefintlig.)"Denna kandidat skulle ge balans till en avdelning som ditt, somredan har så många framstående medlemmar. "(Om du inte redan har en idiot.)"Hans presentation till mitt seminarium förra terminen var verkligen anmärkningsvärt:ett otroligt resultat efter den andra. "(Och vi trodde inte dem heller.)"Hon är helt enhetlig i sin inställning till någon funktion du kan tilldela henne."(I själva verket, till livet i allmänhet ...)
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad de sa:Vad de menade:"Du kommer att ha tur om du kan få honom att arbeta för dig."(Vi säkerligen aldrig lyckats.)Det finns ingen annan anställd som jag kan adekvat jämföra honom.(Jo, våra råttor är inte riktigt anställda ...)"Framgång aldrig kommer att förstöra honom."(Tja, åtminstone inte så mycket mer.)"Man kommer vanligtvis ifrån honom med en bra känsla."(Och en sådan suck av lättnad.)"Hans avhandling är den typ av arbete du förvänta dig inte att se dessa dagar;i det han definitivt har visat sin fullständiga kapacitet. "(Och hans IQ, liksom.)"Han borde gå långt."(Ju längre desto bättre.)"Han kommer att dra full nytta av sin personal."(Han har även en av dem klipper sin gräsmatta efter jobbet.)
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad de säger: Vad de betyder:Ett stort tekniskt genombrott ... Tillbaka till ritbordet.Utvecklad efter år av forskning upptäckte av en ren slump.Projekt bakom ursprungliga tidsplanen på grund Vi arbetar på något annat.oförutsedda svårigheterDesigner är inom tillåtna gränser Vi gjorde det, stretching en punkt eller två.Kundnöjdhet tros Hittills försenat att de ska varaförsäkrade tacksam för någonting alls.Nära samordning projekt Vi ska sprida skulden, campare!Testresultaten var mycket glädjande Det fungerar, och pojke, blev vi förvånade!Designen kommer att slutföras ... Vi har inte börjat ännu, men vi haratt säga något.Hela konceptet har avslagits Killen som konstruerade den sluta.Vi går vidare med ett nytt Vi anlitade tre nya killar, och de ärnärma sparka runt.Ett antal olika metoder ... Vi vet inte vart vi ska, menvi rör oss.Preliminära operativa tester sprängde när vi aktiverat.inconclusiveÄndringar pågår Vi börjar över.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad de säger: Vad de betyder:Nya Olika färger från föregående version.Alla nya Ej kompatibel med tidigare version.Exklusiv Ingen annan har dokumentation.Omatchade Nästan lika bra som tävlingen.Design Enkelhet Företaget skulle inte ge oss några pengar.Idiotsäkert Operation Alla parametrar är hårdkodade.Advanced Design Inget verkligen förstår det.Här äntligen Inte få det gjort i tid.Fält testade vi inte har några simulatorer.År av utveckling Slutligen fick en att arbeta.Oöverträffad prestanda Ingenting någonsin kört långsamt innan.Revolutionerande Disk-enheter att gå runt och runt.Futuristiska körs bara på en nästa generations superdator.Inget underhåll omöjligt att fastställa.Prestanda bevisats arbetat igenom betatestet.Uppfyller tuffa kvalitetsstandarder Det sammanställer utan fel.Garanterad tillfredsställelse Vi skickar dig en annan förpackning om det misslyckas.Lagervara Vi levereras det tidigare och kan göra det igen.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad detta land behöver är en dime som kommer att köpa en bra fem cent bagel.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad detta land behöver är en bra fem cent NÅGOT!
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad detta land behöver är en bra fem cent nickel.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad detta land behöver är en bra fem dollar plasma vapen.
		-- R. Pirsig, "Zen and the Art of Motorcycle Maintenance"

%
Vad vi behöver i detta land, i stället för sommartid, som ingenverkligen förstår i alla fall, är ett nytt koncept som kallas Weekday morgon Time,varvid åtmin 07:00 varje vardag vi går in i ett utrymme lansering-stil "hold" förtvå till tre timmar, under vilken det bara förblir 07:00 På detta sätt kunde vialla vakna upp via en civiliserad gradvis process av stretching och rapningar ochrepor, och det skulle fortfarande vara endast 7:00 när vi var redo att faktisktdyka upp ur sängen.
		-- Dave Barry, "$#$%#^%!^%&@%@!"

%
Vad som inte spikas är min. Vad jag kan bända upp är inte spikas.
		-- Collis P. Huntingdon, railroad tycoon

%
När en Banker hoppar ut genom ett fönster, hoppa efter honom - det är där pengarna finns.
		-- Robespierre

%
När en kollega säger: "Det är inte pengarna utan principen om saken,"det är pengar.
		-- Kim Hubbard

%
När allt annat misslyckas, läs instruktionerna.
		-- Kim Hubbard

%
När jag arbetar, arbetar jag hårt.När jag sitter, sitter jag lätt.Och när jag tänker, går jag sova.
		-- Kim Hubbard

%
När du är osäker, mumla; när de har problem, delegera; när laddning, fundera.
		-- James H. Boren

%
När det inte är nödvändigt att fatta ett beslut, är det nödvändigt att inteta ett beslut.
		-- James H. Boren

%
När rätt sätt, inte semester inte minskar produktiviteten: förvarje vecka du är borta och får ingenting gjort, det finns en annan när din chefär borta och du får dubbelt så mycket gjort.
		-- Daniel B. Luten

%
När chefer prata om att förbättra produktiviteten, de aldrig talarom sig själva.
		-- Daniel B. Luten

%
När lodge mötet bröt upp, Meyer anför till en vän."Abe, jag är i en fruktansvärd knipa Jag är ont om kontanter och jag har inteaning där jag kommer att få det från! ""Jag är glad att höra att" svarade Abe. "Jag var rädd för att dukan ha en uppfattning som du kan låna av mig! "
		-- Daniel B. Luten

%
När du arbetar hårt, få upp och kräkas varje så ofta.
		-- Daniel B. Luten

%
När du inte vet vad de ska göra, gå snabbt och ser orolig.
		-- Daniel B. Luten

%
När du inte vet vad du gör, gör det snyggt.
		-- Daniel B. Luten

%
När du går ut för att köpa, inte visa din silver.
		-- Daniel B. Luten

%
När du gör ditt varumärke i världen, se upp för killar med suddgummin.
		-- The Wall Street Journal

%
När ditt arbete talar för sig själv, inte avbryta.
		-- Henry J. Kaiser

%
Där det finns en vilja finns det en släkting.
		-- Henry J. Kaiser

%
Där det finns en vilja finns det en arvsskatt.
		-- Henry J. Kaiser

%
Även pengar inte kan köpa lycka, låter det verkligen du välja din egenform av elände.
		-- Henry J. Kaiser

%
Även om pengar inte köpa kärlek, uttrycker det du i en stor förhandlingsposition.
		-- Henry J. Kaiser

%
Som utgick ett-lån utgick ett-sörjande.
		-- Thomas Tusser

%
Den som dör med flest leksaker vinner.
		-- Thomas Tusser

%
Varför vara en man när man kan vara en framgång?
		-- Bertolt Brecht

%
Kommer du låna mig $ 20,00 och bara ge mig tio av det?På så sätt kommer du är skyldig mig tio, och jag är skyldig dig tio, och vi kommer att bli ännu!
		-- Bertolt Brecht

%
Önskar utan arbete är som fiske utan bete.
		-- Frank Tyger

%
Arbetet expanderar för att fylla den tillgängliga tiden.
		-- Cyril Northcote Parkinson, "The Economist", 1955

%
Arbetet är av två slag: första, förändra läget för ärendet vid eller närajordytan i förhållande till andra frågor; andra, berätta för andraatt göra så.
		-- Bertrand Russell

%
Arbetet är krabba gräs i gräsmattan i livet.
		-- Schulz

%
Arbeta smartare, inte hårdare, och vara försiktig med din speling.
		-- Schulz

%
Arbete utan en vision är slaveri, är Vision utan arbete en önskedröm,Men vision med arbetet är hoppet om världen.
		-- Schulz

%
XI:Om jorden skulle kunna göras för att rotera dubbelt så fort, chefer skullefå dubbelt så mycket gjort. Om jorden skulle kunna göras för att rotera tjugogånger så snabbt, alla andra skulle få dubbelt så mycket gjort sedan allachefer skulle flyga bort.XII:Det kostar en hel del att bygga dåliga produkter.XIII:Det finns många mycket framgångsrika företag i USA.Det finns också många högavlönade chefer. Policyn är inteblandas de två.XIV:Efter år 2015 kommer det att finnas några flygplanskrascher. Det kommeringa starter heller, eftersom elektronik kommer att uppta 100 procentav varje flygplanets vikt.XV:Den sista 10 procent av prestanda genererar en tredjedel av kostnadenoch två tredjedelar av problemen.
		-- Norman Augustine

%
XLI:Ju mer man producerar, blir mindre ett.XLII:Enkla system är inte möjligt, eftersom de kräver oändlig testning.XLIII:Hårdvara fungerar bäst när det är viktigt att minst.XLIV:Flygplan flygning i 21: a århundradet kommer alltid att vara i en västligriktning, företrädesvis supersonic, korsar tidszoner för att gemertid som behövs för att fastställa trasiga elektronik.XLV:Man bör förvänta sig att den förväntade kan förhindras, menoförutsett skulle ha förväntats.XLVI:En miljard sparas är en miljard intjänas.
		-- Norman Augustine

%
XLVII:Två tredjedelar av jordens yta är täckt med vatten. Den andratredje är täckt med revisorer från huvudkontoret.XLVIII:Ju mer tid du spenderar talar om vad du har gjort, detmindre tid du har att spendera gör vad du har talat om.Så småningom, spenderar du mer och mer tid åt att tala om mindre och mindretills slutligen du lägger all tid åt att tala om ingenting.XLIX:Förordningar växa i samma takt som ogräs.L:Den genomsnittliga reglering har en livslängd en femtedel så länge som enschimpans-talet och en tiondel så länge som en människa - men fyra gångerså länge tjänstemannens som skapade den.LI:Vid tiden för USA Tricentennial, kommer det att finnas merregeringen arbetstagare än det finns arbetare.LII:Personer som arbetar inom den privata sektorn bör försöka spara pengar.Det finns fortfarande möjlighet att det en dag kan vara värdefullt igen.
		-- Norman Augustine

%
XVI:Under år 2054 kommer hela försvarsbudgeten köpa bara enflygplan. Detta flygplan måste delas av flygvapnet ochNavy 3-1 / 2 dagar vardera per vecka med undantag för skottår, när det blirgöras tillgänglig för de flottor för den extra dag.XVII:Mjukvara är som entropi. Det är svårt att förstå, väger ingenting,och lyder termodynamikens andra lag, det vill säga ökar alltid.XVIII:Det är mycket dyrt att uppnå hög opålitlighet. Det är inte ovanligtatt öka kostnaden för ett objekt med en faktor tio för varje faktortio nedbrytning åstadkommes.XIX:Även om de flesta produkter kommer snart att vara för dyrt att köpa, det kommervara en blomstrande marknad för försäljning av böcker om hur man löser dem.XX:Under ett visst år kommer kongressen tillägna den finansieringgodkände föregående år plus tre fjärdedelar av allt ändraadministration förfrågningar - minus 4 procent skatt.
		-- Norman Augustine

%
XXI:Det är lätt att få ett lån om du inte behöver det.XXII:Om aktiemarknaden experter var så expert, skulle de köpa aktier,inte sälja råd.XXIII:Varje uppgift kan fyllas i endast en tredjedel mer tid än vad som ärnärvarande uppskattas.XXIV:Det enda dyrare än stretching schemat för enetablerade projekt accelererar det, som i sig är den mestkostsam åtgärd som människan känner till.XXV:En reviderad tidsplan är att företag vad en ny säsong är att en idrottsmaneller en ny duk till en artist.
		-- Norman Augustine

%
XXVI:Om ett tillräckligt antal hanteringsskikt är överlagrade på varjeandra, kan det säkerställas att katastrofen inte lämnas åt slumpen.XXVII:Rang inte skrämma hårdvara. Inte heller bristen på rang.XXVIII:Det är bättre att vara NYDANARE än reorganizee.XXIX:Chefer som inte producerar framgångsrika resultat håller på att derasjobb bara cirka fem år. De som producerar effektiva resultathänga på ungefär ett halvt decennium.XXX:Vid tiden folk ställer frågorna är redo för svar,de människor som gör arbetet har förlorat kontakten med frågorna.
		-- Norman Augustine

%
XXXI:Den optimala kommitté har inga medlemmar.XXXII:Anställa konsulter för att genomföra undersökningar kan vara ett utmärkt sätt attvrida problem i guld - dina problem i deras guld.XXXIII:Dårar rusa in där etablerade fruktar att beträda.XXXIV:Processen att konkurrens välja entreprenörer att utföra arbetebygger på ett system av belöningar och straff, alla fördeladeslumpmässigt.XXXV:Den svagare tillgängliga uppgifter att grunda en slutsats,desto större noggrannhet som bör citeras för att gedata äkthet.
		-- Norman Augustine

%
XXXVI:Tjockleken på förslag som krävs för att vinna en multimiljonKontraktet är ungefär en millimeter per miljon dollar. Om allaförslag som överensstämmer med denna standard var staplade ovanpå varandralängst ned i Grand Canyon det förmodligen skulle vara en bra idé.XXXVII:Nittio procent av tiden saker blir sämre än förväntat.De övriga 10 procent av den tid du hade rätt att förvänta sig så mycket.XXXVIII:Den tidiga fågeln får masken.Den tidiga mask ... blir uppäten.XXXIX:lovar aldrig att slutföra ett projekt inom sex månader efter utgången avåret - i endera riktningen.XL:De flesta projekten börjar långsamt - och sedan sorts avta.
		-- Norman Augustine

%
Igår var jag en hund. Idag är jag en hund. Imorgon ska jag nog fortfarandevara en hund. Suck! Det finns så lite hopp för avancemang.
		-- Snoopy

%
Du är alltid gör något marginell när chefen droppar av ditt skrivbord.
		-- Snoopy

%
Du kan lura alla människor hela tiden om reklamen är rättoch budgeten är tillräckligt stor.
		-- Joseph E. Levine

%
Du kan berätta för ideal för en nation av dess reklam.
		-- Norman Douglas

%
Du visste jobbet var farligt när du tog den, Fred.
		-- Superchicken

%
Du vet, är skillnaden mellan detta företag och Titanic attTitanic hade betalande kunder.
		-- Superchicken

%
Du eller jag måste ge upp sitt liv till Ahrimanes. Jag skulle hellre det var du.Jag skulle inte tveka att offra mitt eget liv för att skona er, menvi tar lager nästa vecka, och det skulle inte vara rättvist mot företaget.
		-- J. Wellington Wells

%
Du också kan göra stora pengar i den spännande inom pappers SLÄPIG!. Mr Smith Muddla, Mass säger: "Innan jag tog den här kursen jag brukade varaen ödmjuk bitars Twiddler. Nu med vad jag lärde mig på MIT Tech Jag känner verkligenviktig och kan fördunkla och förvirra med det bästa. "Mr Watkins hade följande att säga: "Tio korta dagar sedan allt jag kunde se fram emotatt var en återvändsgränd jobb som ingenjör. Nu Jag har en lovande framtid ochgöra riktigt stora Zorkmids. "MIT Tech kan inte lova dessa fantastiska resultat till alla, men närdu tjänar din MDL examen från MIT Tech din framtid kommer att bli ljusare.SKICKA för vår fria broschyr idag!
		-- J. Wellington Wells

%
