Ditt arbete kommer att fylla en stor del av ditt liv, och det enda sättet att varaverkligen nöjd är att göra vad du tror är stora arbete. Och det enda sättet att görastora arbete är att älska det du gör. Om du inte har hittat det ännu, att se ut.Nöj dig inte. Som med alla frågor av hjärtat, vet du när du hittar den.Och precis som alla bra relation, det bara blir bättre och bättre med årenFortsätt. Så fortsätta leta tills du hittar det. Nöj dig inte.                - Steve Jobs (1955-2011)(1) Undvik stekt kött som arg upp blodet.(2) Om din mage motverkar du, lugna det med häftiga tankar.(3) Håll safter flödar genom klingande runt försiktigt när du flyttar.(4) Gå mycket lätt på laster, såsom att bära på i samhället, somden sociala ramble är inte vilsam.(5) Undvik att köra hela tiden.(6) Do not look back, något kan få på dig.
		-- S. Paige, c. 1951

%
En sammandrabbning av läran är inte en katastrof - det är en möjlighet.
		-- S. Paige, c. 1951

%
Ett moln vet inte varför den rör sig i just en sådan riktning och vid en sådanen hastighet, det känns en impuls ... är detta rätt plats att gå nu. Menhimmel vet orsakerna och mönstren bakom alla moln, och du kommervet också, när du lyfter själv tillräckligt hög för att se bortom horisonter.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
En dröm kommer alltid att segra över verkligheten, när det ges chansen.
		-- Stanislaw Lem

%
En falsk spåman kan tolereras. Men en autentisk soothsayer börskjutas på sikt. Cassandra fick halva sparkar runt hon förtjänade.
		-- R. A. Heinlein

%
Ett stoppat reträttÄr nervpåfrestande och farlig.Att behålla människor som män - och tjänarinnorTar lycka.
		-- R. A. Heinlein

%
En livstid är inte alls tillräckligt länge för att ta reda på vad det handlar om.
		-- R. A. Heinlein

%
Många människor jag känner tror på positivt tänkande, och det gör I. Itro på allt positivt stinker.
		-- Lew Col

%
En man sade till universum:"Sir, finns jag!""Men", svarade universum,"Det faktum inte har skapats i mig en känsla av förpliktelse."
		-- Stephen Crane

%
En befälhavaren ställde frågan: "Vad är vägen?" av ett nyfiket munk."Det är mitt framför ögonen", sade befälhavaren."Varför kan jag inte se det själv?""Eftersom du tänker på dig själv.""Hur du: ser du det?""Så länge du ser dubbelt, säger 'jag inte", och' ni ', och såpå dina ögon är dystra ", sade befälhavaren."När det finns varken 'I' eller 'Du, kan man se det?""När det finns varken 'jag inte heller' Du,som är den som vill se det? "
		-- Stephen Crane

%
En granne kom till Nasrudin, ber att låna hans åsna. "Det är ute pålån "läraren svarade. I det ögonblicket, brayed åsnan högt inutistallet. "Men jag kan höra det Bray, där borta." "Vem tror du"frågade Nasrudin "mig eller en åsna?"
		-- Stephen Crane

%
En präst rådde Voltaire på sin dödsbädd att avstå från djävulen.Svarade Voltaire, "Detta är ingen tid att göra nya fiender."
		-- Stephen Crane

%
En präst frågade: Vad är ödet, Master?Och Mästaren svarade:Det är det som ger en lastdjur sitt existensberättigande.Det är det som män i forna tider var tvungna att bära på ryggen.Det är det som har orsakat länder att bygga stigar från stadenCity på vilka vagnar och bussar passerar, och längs vilken värdshushar kommit att byggas för att avvärja hunger, törst och trötthet.Och det är ödet? sade prästen.Ödet ... Jag tyckte du sa Freight, svarade Mästaren.Det är okej, sade prästen. jag ville vetavad Freight var alltför.
		-- Kehlog Albran, "The Profit"

%
Ett sorgligt spektakel. Om de bebodda, vilken omfattning för misär och dårskap.Om de inte bebodda, vad ett slöseri med utrymme.
		-- Thomas Carlyle, looking at the stars

%
En Scholar frågade sin Mästare, "Mästare, skulle du råda mig om en ordentligkallelse?"Mästaren svarade, "Vissa män kan tjäna sitt hålla med kraften avderas sinnen. Andra måste använda uppgift om deras starka ryggar, ben och händer. Detta ärav samma karaktär som det är med människan. Vissa djur får sin mat lätt,såsom kaniner, svin och getter. Andra djur måste våldsamt kämpar försitt uppehälle, som bäver, mullvadar och myror. Så ni ser, naturkallelse måste passa den enskilde."Men jag har inga förmågor, önskningar, eller fantasi, Mästare", denlärd snyftade.Ifrågasatte mästare ... "Har du tänkt att bli en säljare?"
		-- Thomas Carlyle, looking at the stars

%
En sak är inte nödvändigtvis sant att en människa dör för det.
		-- Oscar Wilde, "The Portrait of Mr. W. H."

%
En blivande lärjunge kom till Nasrudin hydda på berget sida. Menandeatt varje handling av en sådan upplyst är betydande, sökarensåg läraren noga. "Varför du blåser på dina händer?" "Att värmasjälv i kylan. "Senare, Nasrudin hällde skålar varm soppa för sig självoch nykomlingen, och blåste på egen hand. "Varför gör du det, Master?""För att kyla soppan." Det går inte att lita på en man som använder samma processatt komma fram till två olika resultat - varmt och kallt - lärjungen avgick.
		-- Oscar Wilde, "The Portrait of Mr. W. H."

%
Ah, men en mans grepp bör överskrida hans räckhåll,Eller vad är ett himmelrike för?
		-- Robert Browning, "Andrea del Sarto"

%
Alla hoppas överge, ni som skriver här!
		-- Dante Alighieri

%
Alla män vet nyttan av användbara saker;men de vet inte nyttan av meningslöshet.
		-- Chuang-tzu

%
Alla de verkliga saker som jag är på väg att berätta är skamlösa lögner.
		-- The Book of Bokonon / Kurt Vonnegut Jr.

%
Alla vi bör minnas sin orientaliska visdom och hans predikan enZen-liknande avskildhet, som exemplifieras av hans ständiga påminnelse till kontorister,rösträknare, eller andra som växte upphetsad av hans närvaro i sina banker:"Bara ligga ner på golvet och hålla sig lugna."
		-- Robert Wilson, "John Dillinger Died for You"

%
En idé är ett öga från Gud för ser Gud. Vissa av dessa ögonVi kan inte stå ut med att titta ut, vi blinda dem så snabbt som möjligt.
		-- Russell Hoban, "Pilgermann"

%
En idé är inte ansvarig för de människor som tror på den.
		-- Russell Hoban, "Pilgermann"

%
En äldre elev kom till Otis och sa, "Jag har varit att se enstort antal lärare och jag har gett upp ett stort antal nöjen.Jag har fastat varit celibat och stannade vaken nätterna söker upplysning.Jag har gett upp allt jag blev ombedd att ge upp och jag har lidit, menJag har inte upplyst. Vad ska jag göra?"Otis svarade: "Ge upp lidande."
		-- Camden Benares, "Zen Without Zen Masters"

%
Och någonsin har det varit känt att kärlek vet inte sina egna djup tillstimme av separation.
		-- Kahlil Gibran

%
Hur som helst, jag hålla föreställande alla dessa små barn som leker vissa spel i dettastort fält av råg och alla. Tusentals små barn, och ingen är runt -ingen stor, menar jag - utom jag. Och jag står på kanten av någon galenklippa. Vad jag har att göra, jag måste hinna alla om de börjar att gåöver klippan - jag menar om de kör och de ser inte var de ärkommer jag att komma ut från någonstans och fånga dem. Det är allt jag skulle görahela dagen. Jag skulle bara vara Räddaren i nöden. Jag vet det; Jag vet att det är galet,men det är det enda jag skulle verkligen vilja vara. Jag vet att det är galet.
		-- J. D. Salinger, "Catcher in the Rye"

%
Närmar portarna i klostret, Hakuin hittade Ken Zenpredikat till en grupp av lärjungar."Ord ..." Ken orated, "de är men en illusorisk slöja fördunklarden absoluta verklighet - ""Ken!" Hakuin avbrytas. "Din fluga är nere!"Varpå klara ljuset av belysning exploderade på Ken, och hanförångas.På väg till staden, var Hakuin möttes av en ambulerande munk genomsyrasmed andan i morgon."Ah," munken suckade, en saliga leende rynkor över kinderna,"Du är Det ...""Ah", Hakuin svarade pekar ivrigt, "Och Du är fett!"Varpå klara ljuset av belysning exploderade på munken,och han förångas.Därefter sökte guvernören råd Hakuin ropade: "Som vårfiender bär ner på oss, hur skall jag, med en sådan hjärtlös och callowsoldater som jag arvtagare till, hoppas att motstå den överhängande angrepp? ""USA?" snäppas Hakuin.Varpå klara ljuset av belysning exploderade påGuvernör, och han förångas.Sedan gick en redneck upp till Hakuin och förångas den gamla Master medsitt hagelgevär. "Ha! Vispa ya 'till punchline, ya' magra li'l geek!"
		-- J. D. Salinger, "Catcher in the Rye"

%
Arrakis lär attityden hos kniven - hugga av vadofullständig och säger: ". Nu är det fullständig eftersom det slutade här"
		-- Muad'dib, "Dune"

%
Som misslyckanden går, försöker minnas det förflutna är som att försöka greppmeningen med tillvaron. Båda göra en känsla som ett barn klänger påen basket: ens palmer hålla glider.
		-- Joseph Brodsky

%
Vid lågvatten skrev jag en linje på sanden, och gav det hela mitt hjärta och allamin själ. Vid översvämning tidvattnet återvände jag att läsa vad jag hade inskrivet och hittat minokunnighet på stranden.
		-- Kahlil Gibran

%
I slutet av ditt liv det blir en bra vila, och inga ytterligare aktiviteterplaneras.
		-- Kahlil Gibran

%
Vid foten av berget, åska:Bilden av ge näring.den överlägsna mannen är alltså försiktig med sina ordOch tempererade i att äta och dricka.
		-- Kahlil Gibran

%
Skönhet är ett av de sällsynta saker som inte leder till tvivel om Gud.
		-- Jean Anouilh

%
Innan han blev en eremit, var Zarathud en ung präst, ochtog stor glädje i att göra narr av hans motståndare framförhans efterföljare.En dag Zarathud tog sina studenter till en trevlig betesmark ochdär han konfronteras Den sakrala Chao medan hon belåtet bete."Säg mig, du dum odjuret", krävde prästen i hansbefallande röst, "varför inte du göra något värdefullt? Vad är dinSyfte i livet, egentligen? "Mumsa välsmakande gräs, svarade sakrala Chao "MU". (DeKinesiska ideogram för ingen-ting.)När han hörde detta, var absolut ingen upplyst.Främst eftersom ingen förstod kinesiska.
		-- Camden Benares, "Zen Without Zen Masters"

%
Innan du ställa fler frågor, fundera på om du verkligen villveta svaren.
		-- Gene Wolfe, "The Claw of the Conciliator"

%
Brahma sa: Ja, efter att ha hört tio tusen förklaringar, är en dåre intevisare. Men en intelligent man behöver bara två tusen fem hundra.
		-- The Mahabharata

%
Genom protracting liv, vi inte dra ett jota från varaktigheten av döden.
		-- Titus Lucretius Carus

%
Katharsis är något jag förknippar med pornografi och korsord.
		-- Howard Chaykin

%
Visst spelet är riggad.Låt inte det hindra dig; om du inte satsa, kan du inte vinna.
		-- Robert Heinlein, "Time Enough For Love"

%
Chance är kanske Guds verk när han inte ville underteckna.
		-- Anatole France

%
			Kapitel 1Historien hittills:I början universum skapades. Detta har gjort en hel delmänniskor väldigt arga och i stor utsträckning betraktas som ett dåligt drag.
		-- Douglas Adams, HHGG #2, (The Restaurant at the End of the Universe).

%
"Cheshire-Puss", började hon, "vill du berätta för mig, snälla, vilken väg jagborde gå härifrån? ""Det beror en hel del på var du vill komma till", sade katten."Jag bryr mig inte mycket where--" sa Alice."Då spelar det ingen roll vilken väg du går", sade katten.
		-- Douglas Adams, HHGG #2, (The Restaurant at the End of the Universe).

%
Omständigheter härskar män; män utesluter inte omständigheter.
		-- Herodotus

%
Tillfälligheter är andliga vitsar.
		-- G. K. Chesterton

%
Döden är en ande som lämnar en kropp, ungefär som ett skal som lämnar muttern bakom.
		-- Erma Bombeck

%
Döden är Guds sätt att tala om att inte vara en sådan klok kille.
		-- Erma Bombeck

%
Döden är livets sätt att tala om att du har fått sparken.
		-- R. Geis

%
Döden är naturens sätt att återvinna människor.
		-- R. Geis

%
Döden är naturens sätt att säga 'Howdy ".
		-- R. Geis

%
Döden är naturens sätt att tala om att sakta ner.
		-- R. Geis

%
Döden är bara ett sinnestillstånd.Bara den inte lämnar mycket tid att tänka på något annat.
		-- R. Geis

%
Avgår inte från den väg som ödet har tilldelat dig.
		-- R. Geis

%
Beroende på kaninens fot om du vill, men kom ihåg, det hjälpte intekaninen.
		-- R. E. Shay

%
Destiny är en bra sak att acceptera när det går din väg. När det inte är,inte kalla det öde; kalla det orättvisa, förräderi, eller enkel otur.
		-- Joseph Heller, "God Knows"

%
Sjukdom kan botas; öde är obotlig.
		-- Chinese proverb

%
Ditat Deus.[Gud berikar]
		-- Chinese proverb

%
Tror inte på mirakel - lita på dem.
		-- Chinese proverb

%
Misströsta inte av livet. Du har säkert kraft nog för att övervinna dinhinder. Tänk på räven stryker genom trä och fält i en vinternattför något att tillfredsställa sin hunger. Trots kyla och hundar ochfällor, överlever sitt lopp. Jag tror inte någon av dem någonsin begått självmord.
		-- Henry David Thoreau

%
Inte söka döden; död kommer att hitta dig. Men söka den väg som gör dödenen uppfyllelse.
		-- Dag Hammarskjold

%
Ta inte livet för allvarligt; du kommer aldrig att få ut av det levande.
		-- Dag Hammarskjold

%
Gör vad du kan för att förlänga livet, i hopp om att en dag dulära sig vad det är för.
		-- Dag Hammarskjold

%
"Tror du att det finns en Gud?""Jo, ____ någon är ute efter att få mig!"
		-- Calvin and Hobbs

%
Gör din del för att hjälpa till att bevara livet på jorden - genom att försöka bevara din egen.
		-- Calvin and Hobbs

%
Överge inte hopp. Din kapten Midnatt dekoder ring anländer i morgon.
		-- Calvin and Hobbs

%
Överge inte hopp: din Tom Mix dekoder ring anländer i morgon.
		-- Calvin and Hobbs

%
Inte gå till sängs med inget pris på ditt huvud.
		-- Baretta

%
Inte har goda idéer om du inte är villig att vara ansvarig för dem.
		-- Baretta

%
Inte lura dig själv. Lite är relevant, och ingenting varar för evigt.
		-- Baretta

%
Låt inte folk kör du galen när du vet att det är på gångavstånd.
		-- Baretta

%
Gör inte en stor sak av allt; bara ta itu med allt.
		-- Baretta

%
Sluta inte att stampa myror när elefanterna jäktande.
		-- Baretta

%
Ta inte livet på allvar, kommer du aldrig komma ut levande.
		-- Baretta

%
Tvivel är inte motsatsen till tro; Det är en del av tron.
		-- Paul Tillich, German theologian.

%
Ner med kategoriska imperativ!
		-- Paul Tillich, German theologian.

%
På grund av omständigheter utanför din kontroll, är du herre över ditt ödeoch kapten din själ.
		-- Paul Tillich, German theologian.

%
Under resan i livet, kom ihåg att hålla ett öga på en vind i seglen, läktenner under en storm; hagel alla passerande fartyg; och flyga färger stolt.
		-- Paul Tillich, German theologian.

%
Döende är en mycket tråkig, trista angelägenhet. Mitt råd till dig är att hainget som helst att göra med det.
		-- W. Somerset Maugham, his last words

%
Att dö är en av de få saker som kan göras lika lätt liggande.
		-- Woody Allen

%
Varje människa är sin egen fånge i isoleringscell för livet.
		-- Woody Allen

%
Var och en av oss bär sin egen Hell.
		-- Publius Vergilius Maro (Virgil)

%
Antingen jag är död eller min klocka har stannat.
		-- Groucho Marx's last words

%
Även de bästa av vänner inte kan närvara varandras begravning.
		-- Kehlog Albran, "The Profit"

%
Varje människa som nått även hans intellektuella tonåringar börjar misstänkaatt livet är ingen fars; att det inte är elegans komedi ens; att den blommaroch befruktar tvärtom ut ur de djupaste tragiska djupet avväsentlig död i vilken dess motivets rötter försatt. den naturligaarv av alla som är i stånd att andligt liv är en unsubduedskog där varg tjuter och obscena fågel nattchattare.
		-- Henry James Sr., writing to his sons Henry and William

%
Varje person, alla händelser i ditt liv är det att du harlockat dem där. Vad du väljer att göra med dem är upp till dig.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Allt slutar illa. Annars skulle det inte sluta.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Allt i denna bok kan vara fel.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Allt är möjligt. Passera ordet.
		-- Rita Mae Brown, "Six of One"

%
Utför varje handling av thy liv som om det vore din sista.
		-- Marcus Aurelius

%
Expansionsorgan komplexitet; och komplexitet sönderfall.
		-- Marcus Aurelius

%
Fakta är fiende sanningen.
		-- Don Quixote

%
Fain skulle jag klättrar, men fruktar jag att falla.
		-- Sir Walter Raleigh

%
Tro går ut genom fönstret när skönheten kommer in genom dörren.
		-- Sir Walter Raleigh

%
Tron är under vänstra bröstvårtan.
		-- Martin Luther

%
Fyll vad som är tom, tömma det är full, skrapa där det kliar.
		-- Alice Roosevelt Longworth

%
... "Eld" spelar ingen roll, "jord" och "luft" och "vatten" inte spelar någon roll."I" inte spelar någon roll. Inga ord betyder. Men man glömmer verkligheten och minnsord. Ju fler ord han minns, göra smartare sina medmänniskor uppskattar honom.Han ser på de stora omvandlingar av världen, men han ser intedem som de sågs när man såg på verkligheten för första gången.Deras namn kommer till sina läppar och han ler när han smakar dem, tänkte hankänner dem i namngivningen.
		-- Roger Zelazny, "Lord of Light"

%
För snabbverkande lindring, försöka bromsa.
		-- Roger Zelazny, "Lord of Light"

%
För bra, tillbaka bra.Ont, åter rättvisa.
		-- Roger Zelazny, "Lord of Light"

%
För om det är en synd mot liv, består det kanske inte så mycket iförtvivlad av livet som i hopp om ett annat liv och eluding denobevekliga storhet av detta liv.
		-- Albert Camus

%
För din botgöring, säger fem Hail Marys och en högt BLAH!
		-- Albert Camus

%
Force har ingen plats där det finns behov av skicklighet.
		-- Herodotus

%
Fortunes REGLER att leva efter: # 2gås aldrig en järv.
		-- Herodotus

%
FORTUNE regler att leva efter: # 23Skär inte av en polisbil när du gör en olaglig u-sväng.
		-- Herodotus

%
Från att lyssna kommer vishet och från att tala ånger.
		-- Herodotus

%
Från vaggan till kistan underkläder kommer först.
		-- Bertolt Brecht

%
Generellt sett är det långt av krigare beslut acceptans av döden.
		-- Miyamoto Musashi, 1645

%
Att hamna i problem är enkelt.
		-- D. Winkel and F. Prosser

%
Tvillingarna är bara hälften så långt som att få det tillbaka.
		-- D. Winkel and F. Prosser

%
Med tanke på ett val mellan sorg och ingenting, skulle jag välja sorg.
		-- William Faulkner

%
Gud give oss sinnesro att acceptera de saker som vi inte kan förändra, mod attförändra det vi kan, och förstånd att inse skillnaden.
		-- William Faulkner

%
Gud instruerar hjärtat, inte genom idéer, men av smärtor och motsägelser.
		-- De Caussade

%
Gud är tangentpunkten mellan noll och oändligheten.
		-- Alfred Jarry

%
Gud gjorde allt ur ingenting, men intet syns igenom.
		-- Paul Valery

%
Adjö. Jag lämnar eftersom jag är uttråkad.
		-- George Saunders' dying words

%
Adjö, kyler världen.
		-- George Saunders' dying words

%
Fick en ordbok? Jag vill veta meningen med livet.
		-- George Saunders' dying words

%
Stora handlingar består av små handlingar.
		-- Lao Tsu

%
**** Tillväxtcentrum reparationsserviceFör dem som har haft för mycket av Esalen, Topanga, och Kairos. Trött påär äkta hela tiden? Vill du lära dig att vara litefalska igen? Har du avslöjas så mycket att du börjar att undvikapersoner? Har du berört så många människor att de alla börjarkänner detsamma? Gillar att vara lite beroende? Är perfekta orgasmerbörjar tråka ut er? Vill du, för en gångs skull, inte för att uttrycka enkänsla? Eller ännu bättre, inte vara i kontakt med det alls? Kom till oss. Vilovar att befria dig från bördan av din stor potential.
		-- Lao Tsu

%
Lycka är att ha en repa för varje kliar.
		-- Ogden Nash

%
Lycka är bara en illusion, fylld med sorg och förvirring.
		-- Ogden Nash

%
Lycka är att inte ha vad du vill, det vill vad du har.
		-- Ogden Nash

%
Lycka är inte något du upplever; det är något du kommer ihåg.
		-- Oscar Levant

%
Att ha det mest få önskar jag närmast till gudarna.
		-- Socrates

%
Han har visat dig, o människa, vad som är bra. Och vad Herren ber dig,men att göra rättvisa, och att älska vänlighet, och vandrar i ödmjukhet inför din Gud?
		-- Socrates

%
Han är verkligen klokt som vinner visdom från någon annans missöde.
		-- Socrates

%
Han vet inte hur man vet vem vet inte också hur man Okänd.
		-- Sir Richard Burton

%
Han som komponerar själv är klokare än den som komponerar en bok.
		-- B. Franklin

%
Han tänkte på Musashi, Sword Saint, som står i sin trädgård mer äntre hundra år sedan. "Vad är det" Body of a rock '? " Han tillfrågades.Som svar, Musashi kallade en elev av hans och bjuda honom döda sig själv genomslashing hans mage med en kniv. Precis som eleven var på väg att uppfylla,Mästaren stannade handen och sade: "Det är det" Body of a rock "."
		-- Eric Van Lustbader

%
Han som misströstar över en händelse är en fegis, men han som innehar förhoppningar ommänniskans villkor är en dåre.
		-- Albert Camus

%
Den som känner inte och vet att han vet inte är okunnig. Lär honom.Den som känner inte och vet inte att han vet inte är en dåre. Shun honom.Den som känner till och vet inte att han vet sover. Väcka honom.
		-- Albert Camus

%
Han som vet ingenting, vet ingenting.Men den som vet att han vet ingenting vet något.Och den som känner någon vars väns frus bror vet ingenting,han vet något. Eller något sådant.
		-- Albert Camus

%
Han som känner andra är klok.Den som känner sig själv är upplyst.
		-- Lao Tsu

%
Han som vet att enough is enough kommer alltid att ha tillräckligt.
		-- Lao Tsu

%
Den som vet, inte talar. Han som talar, inte vet.
		-- Lao Tsu

%
... Han som skrattar inte tror på vad han skrattar åt, men varkenhan hatar det. Därför skrattar åt det onda inte innebär att förbereda sig förbekämpa den, och skrattar åt bra sätt förneka makt genom vilken bra ärsjälvföröknings.
		-- Umberto Eco, "The Name of the Rose"

%
Här är ett test för att se om ditt uppdrag på jorden är klar:om du lever, är det inte.
		-- Umberto Eco, "The Name of the Rose"

%
Hur kan man bevisa om just nu är vi sover, och alla våratankar är en dröm; eller om vi är vakna, och prata med varandrai vaket tillstånd?
		-- Plato

%
Jag är inte rädd för i morgon, för jag har sett i går och jag älskar idag.
		-- William Allen White

%
Jag trodde inte på reinkarnation i någon av mina andra liv. Jag förstår inte varförJag måste tro på det här.
		-- Strange de Jim

%
Jag vet inte om jag var då en man som drömmer jag var en fjäril, ellerom jag nu en fjäril drömmer jag är en man.
		-- Chuang-tzu

%
Jag söker inte de okunniga; okunniga söka mig - jag kommer att instruera dem.Jag ber bara uppriktighet. Om de kommer ut ur vana, de blir tröttsamt.
		-- I Ching

%
"Jag fick ingenting alls från Supreme upplysningen, och för det mycketAnledningen till att det kallas Supreme upplysningen. "
		-- Gotama Buddha

%
Jag hatar att dö.
		-- Dave Johnson

%
Jag har en enkel filosofi:Fyll vad som är tom.Töm vad är full.Skrapa där det kliar.
		-- A. R. Longworth

%
Jag har ofta ångrat mitt tal, aldrig min tystnad.
		-- Publilius Syrus

%
Jag har sett framtiden och det är precis som den nuvarande, bara längre.
		-- Kehlog Albran, "The Profit"

%
Jag hoppas att du inte låtsas vara ont medan hemlighet är bra.Det skulle vara oärlig.
		-- Kehlog Albran, "The Profit"

%
Jag glömde bara hela mitt livsfilosofi !!!
		-- Kehlog Albran, "The Profit"

%
Jag vet inte hur jag kom in i detta, skall jag kalla det en döende liv eller enlevande död?
		-- St. Augustine

%
"Jag håller helt med dig", sade hertiginnan; "Och den moraliska avdet är - 'Var vad du skulle verkar vara "- eller, om du vill det sättaenklare - `föreställa sig aldrig själv inte att vara annorlunda än vad detkan tyckas andra att vad du var eller kan ha varit var intepå annat sätt än vad du hade skulle varit har dykt upp till dem att varaannat.'"
		-- Lewis Carrol, "Alice in Wonderland"

%
Om en guru faller i skogen med ingen att höra honom, var han verkligen enguru alls?
		-- Strange de Jim, "The Metasexuals"

%
Om en man har en stark tro att han kan njuta av lyxen av skepsis.
		-- Friedrich Nietzsche

%
Om en människa förlorar sin vördnad för någon del av livet, kommer han att förlora sittvördnad för allt liv.
		-- Albert Schweitzer

%
Om jag hade en formel för att kringgå problem, skulle jag inte ge det runt.Problem skapar en förmåga att hantera det. Jag säger inte omfamning problem; det ärlika illa som att behandla det som en fiende. Men jag säger möter den som en vän, fördu se en hel del av det och du hade bättre vara på speaking terms med det.
		-- Oliver Wendell Holmes, Jr.

%
Om jag hade mitt liv att leva över, skulle jag försöka göra fler misstag nästa gång. jagskulle koppla skulle jag limber upp, jag skulle vara dummare än jag har varit härresa. Jag känner väldigt få saker som jag skulle ta på allvar. Jag skulle vara galnare.Jag skulle bestiga fler berg, simma fler floder och titta på fler solnedgångar. jag skulleresa och se. Jag skulle ha fler verkliga bekymmer och färre inbillade.Du förstår, jag är en av dem som bor profylaktiskt och förnuftigtoch förnuftigt, timme efter timme, dag efter dag. Åh, jag har haft mina ögonblick och,om jag hade att göra igen, skulle jag ha mer av dem. I själva verket skulle jag försökerhar ingenting annat. Bara ögonblick, en efter en, i stället för att leva så mångaåren varje dag. Jag har varit en av de människor som aldrig går någonstansutan en termometer, en hotwater flaska, en gurgelvatten, en regnrock och en fallskärm.Om jag hade att göra igen, skulle jag gå platser och göra saker och resorlättare än jag har. Om jag hade mitt liv att leva över, skulle jag börja barfotatidigare på våren och så förbli senare i höst. Jag skulle skolkamer. Jag skulle förmodligen inte göra sådana bra betyg, men jag skulle lära sig mer. jag skullerida på fler merry-go-rundor. Jag skulle plocka fler tusenskönor.
		-- Oliver Wendell Holmes, Jr.

%
Om små gröna män landa i din bakgård, dölja små gröna kvinnordu har i huset.
		-- Mike Harding, "The Armchair Anarchist's Almanac"

%
Om män är inte rädd för att dö,det är till ingen nytta att hota dem med döden.Om män lever i ständig rädsla för att dö,Och om att bryta mot lagen innebär en man kommer att dödas,Vem vågar bryta mot lagen?Det finns alltid en officiell bödel.Om du försöker att ta hans plats,Det är som att försöka vara en mästare snickare och hugga ved.Om du försöker att såga i trä som en mästare snickare,kommer du bara att skada din hand.
		-- Tao Te Ching, "Lao Tsu, #74"

%
Om något ännu inte har gått fel så skulle det i slutändan ha varitfördelaktigt för att det ska gå fel.
		-- Tao Te Ching, "Lao Tsu, #74"

%
Om befälhavaren dör och lärjungen sörjer, liv båda hargått till spillo.
		-- Tao Te Ching, "Lao Tsu, #74"

%
Om sökvägen vara vackra, låt oss inte fråga var den leder.
		-- Anatole France

%
Om det finns en möjlighet till flera saker går fel,den som kommer att orsaka mest skada kommer att vara en att gå fel.Om du uppfattar att det finns fyra möjliga sätt på vilka en procedurkan gå fel, och kringgå dessa, då en femte sätt att snabbt utvecklas.
		-- Anatole France

%
Om det är en synd mot liv, består det kanske inte så mycket i förtvivladav livet som i hopp om ett annat liv och eluding den obevekliga storhetav detta liv.
		-- Albert Camus

%
Om vi ​​inte ändrar vår riktning är vi sannolikt att hamna där vi är på väg.
		-- Albert Camus

%
Om vi ​​inte överleva, behöver vi inte göra något annat.
		-- John Sinclair

%
Om du inte är för dig själv, som kommer att vara för dig?Om du är för dig själv, vad är du?Om inte nu - när?
		-- John Sinclair

%
Om du kan överleva döden, kan du förmodligen överleva någonting.
		-- John Sinclair

%
Om du hittar en lösning och bli fäst vid den, kan lösningen blidin nästa problem.
		-- John Sinclair

%
Om du lura runt med något tillräckligt länge, kommer det så småningom att bryta.
		-- John Sinclair

%
Om du måste hata, hata försiktigt.
		-- John Sinclair

%
Om du måste tänka på det, du har fel.
		-- John Sinclair

%
Om du håller något tillräckligt länge, kan du kasta bort det.
		-- John Sinclair

%
Om du bor tillräckligt länge, kommer du att se att varje seger förvandlas till ett nederlag.
		-- Simone de Beauvoir

%
Om du bara har en hammare, tenderar att se varje problem som en spik.
		-- Maslow

%
Om du skjuta upp det tillräckligt länge, kan det försvinna.
		-- Maslow

%
Om du vägrar att acceptera något annat än det bästa du ofta få det.
		-- Maslow

%
Om du väntar tillräckligt länge, kommer det att gå bort ... efter att ha gjort sin skada.Om det var dåligt, kommer det att vara tillbaka.
		-- Maslow

%
Om du vill ha gudomlig rättvisa, dö.
		-- Nick Seldon

%
Om ditt mål i livet är ingenting, kan du inte missa.
		-- Nick Seldon

%
Om din lycka beror på vad någon annan gör, jag antar att du görhar ett problem.
		-- Richard Bach, "Illusions"

%
Illusionen är den första av alla nöjen.
		-- Voltaire

%
Odödlighet - ett öde värre än döden.
		-- Edgar A. Shoaff

%
I bostad, vara nära marken.I meditation, gräva djupt in i hjärtat.Vid behandling med andra, vara mild och vänlig.I tal, vara sant.I arbetet, vara behörig.I rörelse, vara försiktig med din timing.
		-- Lao Tsu

%
För att upptäcka vem du är, först lära som alla andra är;du vad som finns kvar.
		-- Lao Tsu

%
För att kunna leva fritt och glatt, måste du offra tristess.Det är inte alltid en lätt offer.
		-- Lao Tsu

%
Trots allt, jag tror fortfarande att människor är bra på hjärtat.
		-- Anne Frank

%
I det långa loppet är vi alla döda.
		-- John Maynard Keynes

%
I nästa värld, du är på egen hand.
		-- John Maynard Keynes

%
Faktum är att första ädla sanningen om buddhismen, brukar översättas som`Allt liv är lidande," är mer exakt återges 'liv är fylltmed en känsla av genomträngande otillfredsställelse. "
		-- M. D. Epstein

%
I stället för att älska dina fiender, behandla dina vänner lite bättre.
		-- Edgar W. Howe

%
Intellekt upphäver ödet.Så långt som en människa tänker, är han fri.
		-- Ralph Waldo Emerson

%
Det gör inte att lämna en levande drake av dina beräkningar.
		-- Ralph Waldo Emerson

%
Det är lättare för en kamel för att passera genom ett nålsöga om det ärlätt smord.
		-- Kehlog Albran, "The Profit"

%
Det är Fortune, inte visdom, som styr människans liv.
		-- Kehlog Albran, "The Profit"

%
Det gör inte det vi vill göra, men gillade det vi måste göra,som gör livet välsignade.
		-- Goethe

%
Det är bara genom att riskera våra personer från en timme till en annan att vi leveralls. Och ofta nog vår tro på förhand i en obestyrkt resultatär det enda som gör att resultatet går i uppfyllelse.
		-- William James

%
Det är bara med hjärtat kan man se tydligt; vad som är väsentligt ärosynliga för ögat.
		-- The Fox, 'The Little Prince"

%
Det sägs att den ensamma örnen flyger till bergstoppar medan de ringaant kryper marken, men kan inte själen av myran sväva så högt som örnen?
		-- The Fox, 'The Little Prince"

%
Det är så dum den moderna civilisationen ha gett upp att tro pådjävulen när han är den enda förklaringen till det.
		-- Ronald Knox, "Let Dons Delight"

%
Det är genom symboler som man medvetet eller omedvetet liv och verkoch har sin varelse.
		-- Thomas Carlyle

%
Det kommer att vara fördelaktigt att korsa den stora strömmen ... draken är påvingen på himlen ... den store mannen väcker sig åt sitt arbete.
		-- Thomas Carlyle

%
Det är lättare att ta isär än att sätta ihop det igen.
		-- Washlesky

%
Det är svårt att köra på gränsen, men det är svårare att veta var gränserna går.
		-- Stirling Moss

%
Det är inte verklighet som är viktigt, men hur du uppfattar saker.
		-- Stirling Moss

%
"Det är idag!" sa Nasse."Min favorit dag", sa Puh.
		-- Stirling Moss

%
Det är mycket besvärligt att vara dödlig - du vet aldrig när allt kanplötsligt slutar att hända.
		-- Stirling Moss

%
Joshu: Vad är den sanna vägen?Nansen: Varje sätt är den sanna vägen.J: Kan jag studera det?N: Ju mer du studerar, ju längre från vägen.J: Om jag inte studera det, hur kan jag veta det?N: Vägen tillhör inte saker sett: inte heller saker osynliga.Det hör inte till saker som är kända: eller till saker okända. Dointe söka det, studera det, eller name it. Att hitta dig på den öppnasjälv så bred som himlen.
		-- Stirling Moss

%
Kom bara ihåg, vart du än går, där är du.
		-- Buckaroo Bonzai

%
Vänlighet är början av grymhet.
		-- Muad'dib [Frank Herbert, "Dune"]

%
Låt oss inte se tillbaka i ilska eller framåt i rädsla, men omkring oss i medvetenhet.
		-- James Thurber

%
Livet kan vara så tragiskt - du är här i dag och i morgon.
		-- James Thurber

%
Livet existerar för ingen känd ändamål.
		-- James Thurber

%
Livet är ett stort äventyr - eller det är ingenting.
		-- Helen Keller

%
Livet är att veta hur långt att gå utan passerar linjen.
		-- Helen Keller

%
Livet är som en 10 hastighet cykel. De flesta av oss har växlar vi aldrig använder.
		-- C. Schultz

%
Livet är som en kloak. Vad du får ut av det beror på vad du lagt ned på det.
		-- Tom Lehrer

%
Livet är barndom vår odödlighet.
		-- Goethe

%
Livet är den levande du gör, är död den levande du inte gör.
		-- Joseph Pintauro

%
Livet är lusten att ecstasy.
		-- Joseph Pintauro

%
Livet kan ha någon mening, eller, ännu värre, kan det ha en innebörddu ogillar.
		-- Joseph Pintauro

%
Livet kräver bara från dig den styrka du besitter.Endast en bedrift är möjlig - inte ha rymt.
		-- Dag Hammarskjold

%
Livet suger, men döden inte släcka alls.
		-- Thomas J. Kopp

%
Liksom, om jag inte för mig, då fer shure, som som kommer att vara? Och om du vet,om jag inte gillar fer någon annan, då hej, jag menar, vad är jag? Varom ickenu, som jag vet inte, kanske som när? Och om inte Vem är då jag vet inte, kanskesom Rolling Stones?skrivas Rabbi Hillel.)
		-- Rich Rosen (Rabbi Valiel's paraphrase of famous quote

%
Live aldrig skämmas om något du gör eller säger ärpublicerats runt om i världen - även om vad som publiceras är inte sant.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Att leva i en komplex värld av framtiden är något som att ha binbor i ditt huvud. Men det är de.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Ensamhet är ett fruktansvärt pris att betala för självständighet.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Lång var dagar av smärta jag har tillbringat inom dess väggar, ochlänge var nätterna av ensamhet; och som kan avvika från sinsmärta och hans ensamhet utan ånger?
		-- Kahlil Gibran, "The Prophet"

%
Människans räckvidd överstiga sitt grepp, för varför annars himlen?
		-- Kahlil Gibran, "The Prophet"

%
[Löptid består i upptäckten att] det kommer en kritisk tidpunktdär allt är omvänd, efter vilken punkt blir att förståmer och mer att det är något som inte kan förstås.
		-- S. Kierkegaard

%
Mohandas K. Gandhi ändrade ofta hans sinne offentligt. En medhjälpare en gång frågade honomhur han kunde så fritt motsäga denna vecka vad han hade sagt förra veckan.Den store mannen svarade att det var på grund av denna vecka han visste bättre.
		-- S. Kierkegaard

%
Murphy var en optimist.
		-- Robert Fulghum, "All I ever really needed to know I learned

%
Murphys lag är rekursiv. Tvätta bilen för att göra det regn inte fungerar.
		-- Robert Fulghum, "All I ever really needed to know I learned

%
Musik i själen kan höras av universum.
		-- Lao Tsu

%
Min religion består av en ödmjuk beundran av oändlig överlägsnaande som uppenbarar sig i de små detaljerna vi kan uppfattamed vår bräckliga och svaga sinne.
		-- Albert Einstein

%
Min teologi i korthet är att universum dikterades men inte undertecknat.
		-- Christopher Morley

%
Nasrudin angjort ett stort hus för att samla in för välgörenhet. Tjänaren sade"Min herre är ute." Nasrudin svarade: "Tala om för din mästare att nästa gång hangår ut, bör han inte lämna sitt ansikte i fönstret. Någon kan stjäla den. "
		-- Christopher Morley

%
Nasrudin återvände till sin by från den kejserliga huvudstaden, och bybornasamlades runt för att höra vad som hade passerat. "Vid denna tid," sade Nasrudin, "Jagbara vill säga att kungen talade till mig. "Alla bybor mendummaste sprang för att sprida den underbara nyheter. Den återstående agerfrågade: "Vad gjorde kungen säga till dig?" "Vad han sa - och helt klart,för alla att höra - var "Ut ur min väg!" "The simpleton var överlycklig;Han hade hört ord faktiskt talas av kungen, och sett mycket man detalat med.
		-- Christopher Morley

%
Nasrudin gick in i en butik en dag, och ägaren kom fram för att tjänaHej M. Nasrudin sade, "Först och främst. Såg du mig gå in i ditthandla?"	"Självklart.""Har du någonsin sett mig förut?""Never"."Hur vet du att det var jag?"
		-- Christopher Morley

%
Nasrudin gick in i en tehus och deklamerade, "Månen är mer användbarän solen. ""Varför?", Han frågade."Eftersom på natten vi behöver ljus mer."
		-- Christopher Morley

%
Nasrudin bar hem en bit av levern och receptet för lever paj.Plötsligt en rovfågel svepte ner och ryckte bit kött från hanshand. Som fågeln flög bort, Nasrudin kallas efter det, "dåraktiga fågel! Duhar levern, men vad kan man göra med det utan receptet? "
		-- Christopher Morley

%
Nittio procent av allt är skit.
		-- Theodore Sturgeon

%
Nittio procent av tiden saker bli sämre än du trodde de skulle.De övriga tio procent av den tid du hade rätt att förvänta sig att mycket.
		-- Augustine

%
Ingen människa är en Iland, intire det selfe; varje människa är en peece avKontinent, en del av Maine, om en Clod bi tvättas bort by the Sea,Europa är den lesse, såväl som om en Promontorie var, liksom omen Mannor av dina vänner eller ditt owne var; några bemannar död förminskarmig, eftersom jag är involverad i Mankinde; Och därför aldrig skicka vetaden Klockan klämtar för; Det klämtar för dig.
		-- John Donne, "No Man is an Iland"

%
Vart jag går, är platsen alltid kallat "här".
		-- John Donne, "No Man is an Iland"

%
Ingen användning blir för involverad i livet - du är bara här för en begränsad tid.
		-- John Donne, "No Man is an Iland"

%
Ingen någonsin förstört sin syn genom att titta på den ljusa sidan av något.
		-- John Donne, "No Man is an Iland"

%
Nonsens och skönhet har nära förbindelser.
		-- E. M. Forster

%
Normala tider kan möjligen vara över för alltid.
		-- E. M. Forster

%
Inte varje fråga förtjänar ett svar.
		-- E. M. Forster

%
Ingenting i livet är att frukta. Det är endast för att förstås.
		-- E. M. Forster

%
Ingenting är så enkelt som det verkar vid förstaEller så hopplöst som det verkar i mittenEller som slutade som det verkar i slutändan.
		-- E. M. Forster

%
Ingenting är men det är inte.
		-- E. M. Forster

%
Ingenting är någonsin en total förlust; det kan alltid tjäna som ett dåligt exempel.
		-- E. M. Forster

%
Ingenting är så fast trodde som det som vi stone vet.
		-- Michel de Montaigne

%
Ingenting frågor mycket, och några saker roll alls.
		-- Arthur Balfour

%
Av alla herr elände är bittraste här:att veta så mycket och ha kontroll över ingenting.
		-- Herodotus

%
När tandkrämen är ut ur röret, är det svårt att få det igen.
		-- H. R. Haldeman

%
Väl där bodde en by varelser längs botten av en storCrystal River. Varje varelse i sitt eget sätt höll fast tätt till kvistarnaoch stenar av flodens botten, för att hålla fast var deras sätt att leva, ochmotstå den nuvarande vad varje lärt från födseln. Men en varelsesa till sist, "Jag litar på att den nuvarande vet vart den ska gå. Jag skallsläppa taget och låta det ta mig där det kommer. Klängande, skall jag dö av tristess. "De andra varelser skrattade och sa, "Fool Låt gå, och att den nuvarandedu dyrka kommer att kasta du ramlade och slog över stenarna, och du kommerdör snabbare än tristess! "Men en lyssnade dem inte, och ta ett andetag lät gå, och påen gång ramlade och slog av strömmen över klipporna. Ännu, i tid,som varelsen vägrade att hålla fast igen, lyfte den nuvarande honom fri frånbotten, och han blev slagen och sårad mer.Och varelser nedströms, som han var en främling, ropade, "Seett mirakel! En varelse som själva, men han flyger! Se Messias, komatt rädda oss alla! "Och en transporteras i den aktuella sa," Jag är inte merMessias än du. Floden glädje att lyfta oss fria, om bara vågar vi släppa taget.Vår sanna arbete är denna resa, detta äventyr.Men de ropade mer, "frälsare!" hela tiden klamrar sig faststenar, vilket gör legender av en frälsare.
		-- Richard Bach

%
När du har provat att förändra världen du tycker att det är en massa lättareatt ändra dig.
		-- Richard Bach

%
En dag meddelades att den unge munken Kyogen hade nåtten upplyst tillstånd. Mycket imponerad av denna nyhet, flera av hans kollegorgick för att tala med honom."Vi har hört att du är upplyst. Är detta sant?" hans kollegerstudenter frågade."Det är", svarade Kyogen."Berätta", sa en vän, "hur mår du?""Som eländigt som någonsin", svarade den upplysta Kyogen.
		-- Richard Bach

%
En dag kungen beslutat att han skulle tvinga alla sina undersåtar att berättasanning. En galgen restes framför stadsportarna. En härold meddelade,"Vem skulle komma in i staden måste först svara på sanningen på en frågasom kommer att gå till honom. "Nasrudin var först i kön. Kaptenen påvakt frågade honom: "Vart ska du gå Säg sanningen - den alternativaär döden genom hängning. ""Jag kommer", sade Nasrudin, "att hängas på den galgen.""Jag tror dig inte.""Mycket bra, om jag har ljugit, sedan hänga mig!""Men det skulle göra det sanningen!""Exakt", sade Nasrudin, "din sanning."
		-- Richard Bach

%
Man lär klia där man kan repa.
		-- Ernest Bramah

%
Man möter sitt öde ofta på vägen han tar för att undvika det.
		-- Ernest Bramah

%
En munk sade till den andra, "Fisken har floppat ur nätet! Hur kommer detleva? "Den andra sade," När du har kommit ut ur nätet, ska jag berätta. "
		-- Ernest Bramah

%
Bara att du som är mig kan höra vad jag säger.
		-- Baba Ram Dass

%
Endast de som maklig närma sig som massorna är upptagna påkan vara upptagen om det som massorna ta sköna.
		-- Lao Tsu

%
Paradise är precis som där du är just nu ... bara mycket, mycket bättre.
		-- Laurie Anderson

%
Perfektion uppnås, inte när det inte längre finns något att tillägga, mennär det inte längre finns något att ta bort.
		-- Antoine de Saint-Exupery

%
Kanske den största besvikelser var de du förväntade ändå.
		-- Antoine de Saint-Exupery

%
Filosofi kommer klippa en änglavingar.
		-- John Keats

%
Tryck där den ger och skrapa där det kliar.
		-- John Keats

%
Verkligheten verkar alltid hårdare tidigt på morgonen.
		-- John Keats

%
Verkligheten existerar inte - ännu.
		-- John Keats

%
Verkligheten är illa nog, varför ska jag berätta sanningen?
		-- Patrick Sky

%
Verkligheten är för människor som saknar fantasi.
		-- Patrick Sky

%
Verkligheten är bara en lämpligt mått av komplexitet.
		-- Alvy Ray Smith

%
Verkligheten är bara en krycka för folk som inte kan hantera science fiction.
		-- Alvy Ray Smith

%
Verkligheten är inget annat än en kollektiv föraning.
		-- Lily Tomlin

%
"Verkligheten är den som, när du slutar tro på det, inte försvinner".
		-- Philip K. Dick

%
Kom ihåg, gräshoppa, faller ner 1000 trappan börjar med att snubbla överden första.
		-- Confusion

%
Rule of Life # 1 - Aldrig få skiljas från ditt bagage.
		-- Confusion

%
Se är att tro. Du skulle inte ha sett det om du inte trodde det.
		-- Confusion

%
Eftersom allt i livet är, men en upplevelse perfekt i är vad det är,har ingenting att göra med bra eller dåligt, godtagande eller avvisande, kan man välbrast i skratt.
		-- Long Chen Pa

%
Så lite tid, så lite att göra.
		-- Oscar Levant

%
Ibland även att leva är en handling av mod.
		-- Seneca

%
Ibland får du en nästan oemotståndlig lust att fortsätta leva.
		-- Seneca

%
Standarder är olika för alla ting, så den standard som av människan är avingalunda den enda "säker" standard. Om du förväxla vad som är relativ förnågot säker, har du gått långt från den yttersta sanningen.
		-- Chuang Tzu

%
Lidande ensam existerar ingen som lider;Gärningen finns, men ingen görare därav;Nirvana är, men ingen söker det;Vägen finns, men ingen som reser den.
		-- "Buddhist Symbolism", Symbols and Values

%
Vidskepelse, avgudadyrkan, och hyckleri har gott om löner, men sanningen gåra-tiggeri.
		-- Martin Luther

%
Ta din döende med viss allvar, dock. Skrattar på vägen tilldin utförande är i allmänhet inte förstås av mindre avancerade livsformer,och de kommer att ringa dig galen.
		-- "Messiah's Handbook: Reminders for the Advanced Soul"

%
Att det är är att det inte är är inte.
		-- "Messiah's Handbook: Reminders for the Advanced Soul"

%
Det, det vill säga är.Att det inte är, är det inte.Det, det vill säga är inte det, är det inte.Att det inte är, är inte det, är det.
		-- "Messiah's Handbook: Reminders for the Advanced Soul"

%
Absurda är viktigt begrepp och första sanningen.
		-- A. Camus

%
Det bästa du får är en jämn bryta.
		-- Franklin Adams

%
"Kedjan som kan slet är inte den eviga kedjan."
		-- G. Fitch

%
Den främsta orsaken till problemen är lösningar.
		-- Eric Sevareid

%
Den främsta faran i livet är att du kan ta för många försiktighetsåtgärder.
		-- Alfred Adler

%
Dagarna är tomma och nätterna är overklig.
		-- Alfred Adler

%
Dörren är nyckeln.
		-- Alfred Adler

%
Ögat är ett hot mot fri sikt, är örat ett hot mot subtil hörsel,sinnet är ett hot mot visdom, är varje organ sinnena ett hot mot dessegen kapacitet. ... Fuss, gud Södra oceanen, och Fret, gudeni norra oceanen, hände en gång att träffas i sfären av kaos, gudenom centrum. Chaos behandlade dem mycket vackert och de diskuteras tillsammansvad de kunde göra för att återbetala hans vänlighet. De hade lagt märke till att, medanalla andra hade sju öppningar för syn, hörsel, äta, andas ochså vidare, Chaos hade ingen. Så de bestämde sig för att göra experiment av tråkiga håli honom. Varje dag de borrade ett hål, och på den sjunde dagen dog Chaos.
		-- Chuang Tzu

%
Ju längre du går, desto mindre vet.
		-- Lao Tsu, "Tao Te Ching"

%
Den slutliga vanföreställning är tron ​​att man har förlorat alla illusioner.
		-- Maurice Chapelain, "Main courante"

%
Den första förutsättning för odödlighet är död.
		-- Stanislaw Lem

%
De största sorger är dem vi orsakar oss själva.
		-- Sophocles

%
Den längsta delen av resan sägs vara bortgången av porten.
		-- Marcus Terentius Varro

%
Den stora synd är synd att födas.
		-- Samuel Beckett

%
Märket på din okunnighet är djupet av din tro på orättvisaoch tragedi. Vad larv kallar slutet av världen,mästare kallar en fjäril.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Ju fler lagar och ordning görs framträdande, desto fler tjuvar ochrånare kommer det att finnas.
		-- Lao Tsu

%
Ju mer du klaga, låter längre Gud du bor.
		-- Lao Tsu

%
Mossan på trädet inte frukta klor av Hawk.
		-- Lao Tsu

%
Den mest kostsamma av alla galenskaper är att tro passionerat i påtagligtinte sant. Det är den högsta ockupationen av mänskligheten.
		-- H. L. Mencken

%
Den enda skillnaden mellan en brunst och en grav är deras dimensioner.
		-- H. L. Mencken

%
Den enda lycka ligger i anledning; resten av världen är dyster.Den högsta orsaken, men jag ser i arbete konstnär, och han kanuppleva det som sådant. Lycka ligger i snabbhet känsla ochtänker: resten av världen är långsam, gradvis och dum. Vem som änkunde känna loppet av en ljusstråle skulle bli mycket glad, för det är mycketsnabb. Att se sig själv ger lite glädje. Om däremot känns enmycket glädje i detta, är det på grund på botten man inte tänker påsjälv men av ett ideal. Detta är långt, och endast snabba skall nådet och är glada.
		-- Nietzsche

%
Optimisten tror att detta är den bästa av alla tänkbara världar,och pessimisten vet det.
		-- J. Robert Oppenheimer, "Bulletin of Atomic Scientists"

%
Ändå bekännelser menar mycket lite, coth svarade mörka gud, ännu taladenästan försiktigt. Optimisten proklamerar att vi lever i den bästa av allavärldar; och pessimisten fruktar att detta är sant.
		-- James Cabell, "The Silver Stallion"

%
Dikterna, alla tre hundra av dem, kan sammanfattas i en av sina fraser:"Låt våra tankar vara korrekt".
		-- Confucius

%
Priset för framgång i filosofi är trivialitet.
		-- C. Glymour.

%
Frågorna förblir desamma. Svaren är evigt variabel.
		-- C. Glymour.

%
Loppet är inte alltid den snabba, eller kampen för att den starka, mendet är så att satsa.
		-- Damon Runyon

%
Roten till allt vidskepelse är att män observera när en sak träffar,men inte när det missar.
		-- Francis Bacon

%
Frälsaren blir offer.
		-- Francis Bacon

%
Själen skulle ha någon regnbåge hade ögonen inga tårar.
		-- Francis Bacon

%
Tillståndet för oskuld innehåller bakterier av alla framtida synd.
		-- Alexandre Arnoux, "Etudes et caprices"

%
Den sanna vägen går över ett rep som inte är sträckt vid någon hög höjdmen strax ovanför marken. Det verkar mer för att göra folk snubblarän att beträdas.
		-- Franz Kafka

%
Sanningen är sällan ren och aldrig enkel.
		-- Oscar Wilde

%
Sanningen är vad är; vad som borde vara är en smutsig lögn.
		-- Lenny Bruce

%
Sanningen om en sak är känslan av det, inte tänka på det.
		-- Stanley Kubrick

%
Sanningen du talar har inget förflutet och ingen framtid. Det är, och det är allt detbehöver vara.
		-- Stanley Kubrick

%
Världen är din motion-bok, de sidor där du gör dina summor.Det är inte verkligheten, även om du kan uttrycka verkligheten finns om du vill.Du är också fri att skriva nonsens eller lögner, eller att riva sidorna.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Det finns inga som helst olyckor i universum.
		-- Baba Ram Dass

%
Det finns inga vinnare i livet, enda överlevande.
		-- Baba Ram Dass

%
Det finns tio eller tjugo grundläggande sanningar, och livet är en process förupptäcka dem om och om och om igen.
		-- David Nichols

%
Det finns mer i livet än att utöka dess hastighet.
		-- Mahatma Gandhi

%
Det finns ingen tröst utan smärta; sålunda definierar vi frälsning genom lidande.
		-- Cato

%
Det finns inget botemedel mot födelse och annat än att njuta av intervallet död.
		-- George Santayana

%
Det finns ingen synd, men okunnighet.
		-- Christopher Marlowe

%
Det finns inget som inte kan besvaras med hjälp av min lära ", sägeren munk, som kommer in i ett tehus där Nasrudin satt."Och ändå bara en kort tid sedan, jag utmanades av en lärd medett ovedersägligt fråga ", säger Nasrudin."Jag kunde ha svarat det om jag hade varit där.""Mycket bra. Han frågade:" Varför är du bryta sig in i mitt hus imitt i natten? "
		-- Christopher Marlowe

%
Det finns bara ett allt.
		-- Christopher Marlowe

%
Att få något rent, måste man få något smutsigt.Att få något smutsigt, behöver man inte att få något ren.
		-- Christopher Marlowe

%
Att ge lycka är att förtjäna lycka.
		-- Christopher Marlowe

%
Att ge av sig själv, måste du först känna dig själv.
		-- Christopher Marlowe

%
Ha dött en gång är tillräckligt.
		-- Publius Vergilius Maro (Virgil)

%
Att leda människor, måste du följa bakom.
		-- Lao Tsu

%
Sanning inte har någon särskild tid för sig. Dess timme är nu - alltid.
		-- Albert Schweitzer

%
Sanningen är svårt att hitta och svårare att oklar.
		-- Albert Schweitzer

%
Sanningen aldrig kommer till världen men som en oäkting, till smälekav honom som förde hennes födelse.
		-- Milton

%
Två män kom innan Nasrudin när han var domare. Den första mannen sa,"Den här mannen har bitit mitt öra - Jag kräver ersättning." Den andra mannen sa,"Han bet det själv." Nasrudin drog sig tillbaka till sina kammare, och tillbringade en timmeförsöker bita hans eget öra. Han lyckades bara välter och blåmärkenpannan. Återvänder till rättssalen, uttalas Nasrudin, "Undersökman vars öra blev biten. Om pannan blåmärken, gjorde han det själv ochfallet avslås. Om pannan inte är skadade, gjorde den andre detoch måste betala tre silver bitar. "
		-- Milton

%
Två män satt över kaffe, överväger vilken typ av saker,med all respekt för deras frukost. "Jag undrar varför det är atttoast alltid faller på smörade sidan ", sade en."Säg mig", svarade hans vän, "varför du säger en sådan sak. Tittapå detta. "Och han tappade sin skål på golvet, där det landade påtorra sidan."Så, vad har du att säga till din teori nu?""Vad ska jag säga? Du smörad uppenbarligen fel sida."
		-- Milton

%
Avfall inte färska tårar över gamla sorger.
		-- Euripides

%
Vi kan förkroppsliga sanningen, men vi kan inte veta det.
		-- Yates

%
Vi har ingen annanstans att gå ... detta är allt vi har.
		-- Margaret Mead

%
Vi har bara två saker att oroa sig: Att det aldrig kommer att fåtillbaka till det normala, och att de redan har.
		-- Margaret Mead

%
Vi har anledning att vara rädd. Detta är en fruktansvärd plats.
		-- John Berryman

%
Vi finner sällan någon som kan säga att han har levt ett lyckligt liv, och sominnehåll med sitt liv, kan gå i pension från världen som en nöjd gäst.
		-- Quintus Horatius Flaccus (Horace)

%
Vi är alla i detta ensam.
		-- Lily Tomlin

%
Vi är dödliga - det vill säga, vi är okunniga, dumma, och syndig -men de är bara nackdelar. Vår stolthet är att ändå nu ochdå, vi gör vårt bästa. Ett par gånger vi lyckas. Vad mer vågar vi begära?
		-- Ensign Flandry

%
"Vi pratar inte om samma sak", sade han. "För dig världen ärkonstigt eftersom om du inte är uttråkad med det du är på kant med det. För migvärlden är konstigt eftersom det är häpnadsväckande, enormt, mystisk,outgrundlig; mitt intresse har varit att övertyga dig om att du måste accepteraansvar för att vara här, i denna fantastiska värld, i denna fantastiskaöken, i denna underbara tid. Jag ville övertyga dig om att du måstelära sig att göra varje handling räknas, eftersom du kommer att vara här för endast enkort stund, i själva verket, för kort för att bevittna alla underverk det. "
		-- Don Juan

%
Tja, tänkte han, eftersom varken aristoteliska Logic eller disciplinernaof Science tycktes erbjuda mycket hopp, är det dags att gå bortom dem ...Dra några djupa jämna andetag, gick han ett mentalt tillstånd praktiserasendast av Masters of the Universal Way of Zen. I det hans sinne flöt fritt,kunna rota efter behag bland bitar av data som han hade absorberats,ostörd av någon yttre störningar. Logiska strukturer inte längrehämmade honom. Pre-föreställningar, fördomar, försvann vanliga mänskliga normer.Allt, de tidigare trivialt liksom de en gång trodde viktig,blev helt lika genom att förvärva ett absolut värde, avslöjar relationerinte uppenbart för vanlig syn. Som pärlor uppträdda på ett snöre av sina egnamening, pekade varje sak till sin egen utrett av tillvaron, som delas avalla. Slutligen, varje började smälta i varje, bor själv samtidigt som de bliralla andra. Och Sinne inte längre övervägs problem, men blev problem,förstöra subjekt-objekt genom att bli dem.Tiden gick, obeaktade.Slutligen, fanns det en trevande omröring, varefter en avgörande en, ochNakamura uppstod ett leende på läpparna och mot bakgrund av skratt i hans ögon.
		-- Wayfarer

%
Tja, du vet, oavsett var du går, där är du.
		-- Buckaroo Banzai

%
"Jo", Brahma sa, "även efter tio tusen förklaringar, är en dåre inteklokare, men en intelligent man kräver endast två tusen fem hundra. "
		-- The Mahabharata.

%
Vad inte förstör mig, gör mig starkare.
		-- Nietzsche

%
Vad gör universum så svårt att förstå är att det finns ingetatt jämföra den med.
		-- Nietzsche

%
Vad vettig människa kan leva i den här världen och inte vara galen?
		-- Ursula K. LeGuin

%
Vad vi är Guds gåva till oss.Vad vi Bli är vår gåva till Gud.
		-- Ursula K. LeGuin

%
Oavsett sker från kärlek är alltid bortom gott och ont.
		-- Friedrich Nietzsche

%
Oavsett vad du gör kommer att vara obetydlig, men det är mycket viktigt att du gör det.
		-- Gandhi

%
När det är mörkt nog kan du se stjärnorna.
		-- Ralph Waldo Emerson,

%
När högtalaren och han vem han är talar inte förstår, är attmetafysik.
		-- Voltaire

%
När vinden är stor, båge innan den;när vinden är tung, ge efter för det.
		-- Voltaire

%
När du är ung, du njuta av en ihållande illusion som förr eller senarenågot fantastiskt kommer att hända, att ni kommer att överskridadina föräldrars begränsningar ... Samtidigt känner du säker på att det i allaöknen möjlighet; i alla skogar åsikt, det finns envital något som kan vara känd - kända och gripas. Att vi kommersmåningom vet det, och konvertera hela mysteriet till en sammanhängandeberättelse. Så att då en sanna liv - den punkt på allt -kommer att dyka upp från dimman i ett rent ljus, i total förståelse.Men det är inte som att alls. Men om det inte är, där kom idénfrån att tortera och oroa oss?
		-- Brian Aldiss, "Helliconia Summer"

%
När du dör, förlorar du en mycket viktig del av ditt liv.
		-- Brooke Shields

%
Som inte litar tillräckligt kommer inte att lita på.
		-- Lao Tsu

%
Visdom är att veta vad man ska göra med vad du vet.
		-- J. Winter Smith

%
Visdom är sällan på bästsäljarlistan.
		-- J. Winter Smith

%
[Visdom] är en livets träd för dem omtag i henne, gör gärna vart och ett håller henne snabbt.
		-- Proverbs 3:18, NSV

%
Med lyssna kommer vishet, med talande ånger.
		-- Proverbs 3:18, NSV

%
Wonder är känslan av en filosof, och filosofi börjar i under.[Va? Det är som Johnson citerar Boswell]
		-- Socrates, quoting Plato

%
	Jobba hårt.	Rocka hårt.Ät hårt.Sömn Hård.Grow Big.Glasögon om du behöver 'Em.
		-- The Webb Wilder Credo

%
Ja, men som själv vill du vara?
		-- The Webb Wilder Credo

%
Du aldrig gett en önskan utan också med tanke på denmakt att göra det är sant. Du kanske måste arbeta för det, dock.Advanced Soul "
		-- R. Bach, "Messiah's Handbook : Reminders for

%
Du kan alltid plocka upp din nål och flytta till en annan spår.
		-- Tim Leary

%
Du kan få * någonstans * i tio minuter om du kör tillräckligt snabbt.
		-- Tim Leary

%
Du kan aldrig tala om vilken väg tåget gick genom att titta på spåren.
		-- Tim Leary

%
Du kan inte längre vinna ett krig än du kan vinna en jordbävning.
		-- Jeannette Rankin

%
Du kan observera en hel del bara genom att titta på.
		-- Yogi Berra

%
Du kan bara leva en gång, men om du gör det rätt, är en gång tillräckligt.
		-- Yogi Berra

%
Du kan inte komma dit härifrån.
		-- Yogi Berra

%
Du kan inte laga en armbandsur medan faller från ett flygplan.
		-- Yogi Berra

%
Du kan inte trycka på en sträng.
		-- Yogi Berra

%
Du kan inte springa iväg för evigt,Men det är inget fel med att få en bra försprång.
		-- Jim Steinman, "Rock and Roll Dreams Come Through"

%
"Du kan inte överleva genom att suga saften från en våt vante."		   Om och om igen"
		-- Charles Schulz, "Things I've Had to Learn Over and

%
Du kan inte ta den med dig - särskilt när de passerar en statsgränsen.
		-- Charles Schulz, "Things I've Had to Learn Over and

%
Du klättra för att nå toppen, men när det upptäcker att alla vägarleder ner.
		-- Stanislaw Lem, "The Cyberiad"

%
Du har all evighet att vara försiktig med när du är död.
		-- Lois Platford

%
Du måste köra så fort du kan bara stanna där du är.Om du vill komma någonstans, måste du springa mycket snabbare.
		-- Lewis Carroll

%
"Du menar, om du tillåter befälhavaren att vara ohövlig, att behandla dignågot gammalt sätt han vill, och att förolämpa din värdighet, då han finner digpassar att höra hans syn på saken? ""Tvärtom. Du måste försvara din integritet, förutsattdu har integritet att försvara. Men du måste försvara den ädelt, inte avimitera sin egen låg beteende. Om du är försiktig när han är grov,om du är artiga där han är ouppfostrad, då han kommer att känna igen dig sompotentiellt värda. Om han inte gör det, då är han inte en mästare, trots allt,och du kan gärna spöa honom. "
		-- Tom Robbins, "Jitterbug Perfume"

%
Du kommer alltid att hitta något i den sista platsen du ser ut.
		-- Tom Robbins, "Jitterbug Perfume"

%
"Du skulle göra klokt i att inte föreställa sig djup", sade han. "Allt som verkarav viktig händelse bör bodde på som om det var av liten anmärkning.Omvänt måste trivialiteter skötas med största omsorg.Eftersom döden är betydelsefull, ge det ingen tanke; eftersom seger är viktig,ge det ingen tanke; eftersom metoden av prestation och upptäckt är mindrebetydelsefulla än effekten, uppehållstid alltid på metoden. Du kommer att stärkasjälv på det här sättet. "
		-- Jessica Salmonson, "The Swordswoman"

%
Din lycka är sammanflätad med din syn på livet.
		-- Jessica Salmonson, "The Swordswoman"

%
Ditt sinne förstår vad du har lärt; ditt hjärta, vad som är sant.
		-- Jessica Salmonson, "The Swordswoman"

%
Din enda skyldighet i någon livstid är att vara sann mot dig själv. Varelsesant till någon annan eller något annat är inte bara omöjligt, men dettecken på en falsk messias. De enklaste frågorna är de mest djupgående.Var föddes du? Var är ditt hem? Vart är du på väg? Vadgör du? Tänk på dessa en gång i en stund och titta på dina svarändra.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Din bild av världen förändras ofta precis innan du får den i fokus.
		-- Messiah's Handbook : Reminders for the Advanced Soul

%
Din peruk styr spelningen.
		-- Lord Buckley

%
Du kan marschera till takten av en annan trummis, men du ärfortfarande i paraden.
		-- Lord Buckley

%
Universum består av berättelser, inte av atomer.
		-- Muriel Rukeyser

%
Frihet är vad du gör med vad som gjorts för dig.
		-- Jean-Paul Sartre

%
Det finns en hemlig person som oskadad inom varje individ.
		-- Paul Shepard

%
Vi styrs inte av arméer och polisen men av idéer.
		-- Mona Caird, 1892

%
Den första regeln för alla intelligenta mixtrande är att hålla alla delar.
		-- Aldo Leopold, quoted in Donald Wurster's "Nature's Economy"

%
Du måste vara ändringen som du önskar att se i världen.
		-- Mahatma Gandhi

%
Inga människor är dåliga, precis som ingen är allt bra.Tecumseh, (Shawnee) till sin brorson Spemica Lawba 1790
		-- Mahatma Gandhi

%
Min anledning säger att mark kan inte säljas - ingenting kan säljas utansådant som kan transporteras bort. Black Hawk (Saulk)
		-- Mahatma Gandhi

%
Sälja ett land! Varför inte sälja luften, det stora havet, liksomjord? Inte den store Anden göra dem alla för att använda hansbarn? Tecumseh, (Shawnee)
		-- Mahatma Gandhi

%
Befria dig från negativ påverkan. Negativa tankar är gamlavanor som gnaga på rötterna av själen.Moses Shongo, (Seneca)
		-- Mahatma Gandhi

%
... Allt på denna jord har ett syfte, varje sjukdom en ört att botadet, och varje människa ett uppdrag. Detta är den indiska teorin om tillvaron.Sörjande duva, (Salish 1888-1936)
		-- Mahatma Gandhi

%
"Der bestirnte Himmel über mir und das moralische Gesetz i mir"det är"Den stjärnhimlen ovanför mig, och den moraliska lagen i mig."
		-- The epigraph on Kant's tombstone.

%
Orden flyga iväg, skrifter kvar.
		-- The epigraph on Kant's tombstone.

%
Jag är vad du kommer att vara; Jag var vad du är.
		-- The epigraph on Kant's tombstone.

%
Folket härskar.
		-- The epigraph on Kant's tombstone.

%
Kanske minnet av dessa saker kommer att visa en källa till framtidanöje.
		-- Virgil

%
Någon som förstår allt som kommer ut ur förmögenhet förmodligenhar ett problem
		-- Virgil

%
Om en miljon människor säger en dum sak, är det fortfarande en dum sak.
		-- Anatole France

%
"Få synder är mindre förlåtligt i artigt samhället än att erbjuda dålig folk produkter de aktivt söker. "   - Katherine Mangu-Ward, "Utbildning för vinst", Reason Magazine, juli 2008
		-- Anatole France

%
Din tid är begränsad, så slösa inte det levande någon annans liv                - Steve Jobs (1955-2011)
		-- Anatole France

%
