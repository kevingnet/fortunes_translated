En bok är ett verk av ett sinne, gör sitt arbete på det sätt som ett sinne anserbäst. Det är farligt. Är ett verk av några enbart individuella sinne sannolikttjäna syftena med kollektivt accepterade kompromisser, som är kända inomskolor som "standarder"? Alla ihåg att audaciously skulle sätta sig tillbaka tillarbeta ensam är säkert ett dåligt exempel för eleverna, och förmodligen, ominte rent antisocial, åtminstone en lite utanför centrum, självsvåldiga,elitistisk. ... Det är bara bra pedagogik, därför att hålla sig borta från sådanasaker, och användning i stället, om filmremsor och rap-sessioner måste varakompletteras "texter" väljs eller framställas, eller anpassas, genom verkligproffs. Dessa texter kallas "läsning". De är deakademiska motsvarigheten till "lyssnande material" som fyller väntsalar,och "äta material" som du kan köpa i tusentals bekvämt ätaresurscentra längs vägarna.
		-- The Underground Grammarian

%
En definition av undervisningen: gjutning falska pärlor för riktiga svin.
		-- Bill Cain, "Stand Up Tragedy"

%
En dåre hjärna smälter filosofi i galenskap, vetenskap i vidskepelse, ochkonst i pedanteri. Därför Högskoleutbildning.
		-- G. B. Shaw

%
En bra fråga är aldrig besvarad. Det är inte en bult som skall dras åtpå plats men ett frö att planteras och bära mer frö mothopp om grönare landskap idé.
		-- John Ciardi

%
En grammatiker liv är alltid i spänd.
		-- John Ciardi

%
Ett stort antal människor tror att de tänker när de är baraordna sina fördomar.
		-- William James

%
En mamma mus tog sin stora kull för en promenad över köketvåning en dag när den lokala katten, genom en bedrift av stealth ovanlig även fördess art, lyckats fånga dem i ett hörn. Barnen kröp,livrädd av denna skräckinjagande besten, klagande gråt, "Hjälp, mor!Rädda oss! Rädda oss! Vi är rädda, mor! "Mor mus, med den hopplösa tapperhet en förälder skydda sinbarn, vände med tänderna blottade till katten, tornar enorma ovanför dem,och plötsligt började skälla på ett sätt som skulle ha gjort någon Dobermanstolt. Den överraskad katt flydde i skräck för sitt liv.Som hennes tacksam avkomma flockades runt hennes skrika "Åh, mamma,du räddade oss! "och" Yay! Du skrämde katten away! "Vände hon sig till demmålmedvetet och sade: "Du ser hur bra det är att känna en andraspråk?"
		-- William James

%
En liknelse of Modern forskning:Bob har förlorat sina nycklar i ett rum som är mörk med undantag för enupplysta hörn."Varför ser du under ljuset, du tappade dem i mörkret!""Jag kan bara se här."
		-- William James

%
En penna med någon punkt behöver ingen suddgummi.
		-- William James

%
En plan för förbättring av engelska stavningskrivs Mark TwainTill exempel, i år en som värdelös bokstaven "C" skulle tas bortsom skall replased antingen med "k" eller "s", och på samma sätt "x" skulle inte längrevara en del av alfabetet. Den enda Kase där "c" skulle behållasskulle vara den "ch" formation, som kommer att behandlas senare. år 2kan reformera "w" stavning, så att "som" och "en" skulle tasamma konsonant, LIST År 3 kan mycket väl avskaffa "y" replasing det med"I" och Iear 4 kanske fiks den "g / j" anomali wonse för alla.Jenerally, då skulle förbättringen kontinue iear bai iearmed Iear 5 gör awai med onödiga dubbla konsonants och Iears 6-12eller så modifaiing vowlz och rimeining voist och unvoist konsonants.Bai Iear 15 eller sou, wud det fainali bi posibl tu Meik ius ov thiridandant letez "c", "y" och "x" - bai nu Jast en Memori i maindzov Ould doderez - tu riplais "ch", "sh", och "th" rispektivli.Fainali, xen, aafte sam 20 IERS ov orxogrefkl riform, wi Wudhev en lojikl, werld kohirnt speling i ius xrewawt xe Ingliy-spiking.
		-- William James

%
En professor är den som talar i någon annans sömn.
		-- William James

%
En läsare rapporterar att när patienten dog, den behandlande läkarenregistreras följande på patientjournalen: "Patient underlåtit att uppfyllahans välbefinnande potential. "En annan läkare rapporterar att i ett färskt nummer av den * American Journalof Family Practice * loppor kallades "blodsugande leddjur vektorer."En läsare rapporterar att armén kallar dem "vertikalt utplacerade anti-personal enheter. "Du kallar dem förmodligen bomber.På McClellan Air Force bas i Sacramento, Kalifornien, civilmekanik placerades på "icke-duty, icke-pay status." Det vill säga, de sparken.Efter att ha tagit resan under en livstid, skickade våra läsare hans tolv rullarfilm till Kodak för att utveckla (eller "behandling", som Kodak gillar att kalla det)bara för att få följande meddelande: "Vi måste konstatera att under hanteringenav dina tolv 35mm Kodachrome glid order, var filmerna inblandade i enovanlig laborativ erfarenhet. "Användningen av den passiva är en särskilt trevligberöring, tycker du inte? Ingen gjorde något till filmerna; de hade bara en dåligerfarenhet. Naturligtvis våra läsare kan alltid gå tillbaka till Tibet och ta hansbilder på nytt med hjälp av tolv ersättare rullar Kodak så generöstsänt honom.
		-- Quarterly Review of Doublespeak (NCTE)

%
En student som ändrar historiens förmodligen tar en examen.
		-- Quarterly Review of Doublespeak (NCTE)

%
En synonym är ett ord som du använder när du inte kan stava det ord du försttänkte på.
		-- Burt Bacharach

%
En tautologi är en sak som är tautologier.
		-- Burt Bacharach

%
Ett universitet är vad en högskola blir då fakulteten tappar intressethos eleverna.
		-- John Ciardi

%
"En universitet utan studenter är som en salva utan en fluga."
		-- Ed Nather, professor of astronomy at UT Austin

%
Om alla vissa män åstadkomma i livet är att skicka en son till Harvard.
		-- Ed Nather, professor of astronomy at UT Austin

%
Abstrakt:Denna studie undersökte förekomsten av slips täthet mellan en gruppav 94 vita kragen arbetande män och effekten av en tät affärs skjortkrageoch slips på det visuella resultatet för 22 manliga försökspersoner. Av tjänstemänmän mäts var 67% befunnits vara klädd slips som var hårdare änhalsen omkrets. Den visuella diskriminering av de 22 försökspersoner varutvärderas med hjälp av en testfrekvens kritisk flimmer (CFF). Resultaten av CFFtestet indikerade att snäva slips minskat betydligt den visuellaprestanda av de ämnen och att visuella prestanda inte förbättraomedelbart när tight slips avlägsnades.Hals i förhållande till Visual Performance. "Human Factors 29,# 1 (februari 1987), pp. 67-71.
		-- Langan, L. M. and Watkins, S. M. "Pressure of Menswear on the

%
Akademiska politik är den mest onda och bittra form av politik,eftersom insatserna är så låg.
		-- Wallace Sayre

%
Akademiker vård, det är som.
		-- Wallace Sayre

%
=============== ALLA FRESHMEN OBS ===============För att minimera schemaläggning förvirring, vänligen inse att om du tar enkurs som erbjuds endast en gång på en viss dag, och en annan som ärerbjuds på alla gånger på samma dag, kommer den andra klassen ordnas som tillråd maximal olägenhet för studenten. Till exempel, om du råkaratt arbeta på campus, kommer du att ha 1-2 timmar mellan klasser. Om du pendlar,kommer det att finnas minst 6 timmar mellan de två klasserna.
		-- Wallace Sayre

%
En investering i kunskap betalar alltid det bästa intresse.
		-- Benjamin Franklin

%
Eventuella två filosofer kan berätta för varandra allt de har två timmar.
		-- Oliver Wendell Holmes, Jr.

%
Som general de Gaulle erkänner occassionally Amerika att vara dotterEuropa, så jag är glad att komma till Yale, dotter till Harvard.
		-- J. F. Kennedy

%
Så länge som svaret är rätt, vem bryr sig om frågan är fel?
		-- J. F. Kennedy

%
I korthet resultaten är att när du presenteras med en raddata- eller en sekvens av händelser i vilka de instrueras att upptäckaen underliggande order, ämnen visar starka tendenser att uppfatta ordningoch kausalitet i slumpmässiga matriser, för att uppfatta ett mönster eller korrelationsom verkar a priori intuitivt korrekt även när den faktiska korrelationeni data är bakvända, att dra förhastade slutsatser om rätthypotes, att söka och använda endast positiva eller bekräftande bevis förtolka bevis frikostigt som bekräftande, misslyckas med att generera ellerutvärdera alternativa hypoteser, och har därmed lyckats att utsätta sigendast bekräftande fall vara falskeligen utge säker på giltighetenav sina domar (Jahoda, 1969; Einhorn och Hogarth, 1978). ianalys av tidigare händelser, är dessa tendenser förvärras av bristandeuppskatta fallgropar post hoc-analyser.
		-- A. Benjamin

%
Brittisk utbildning är förmodligen den bästa i världen, om du kan överlevaDet. Om du kan inte det finns någonting kvar för dig men den diplomatiska kåren.
		-- Peter Ustinov

%
... Men om vi skrattar med hån, vi kommer aldrig att förstå. Mänskligintellektuell kapacitet har inte ändrats i tusentals år, eftersomvi kan berätta. Om intelligenta människor investerat intensiv energi i frågorsom nu verkar dumt för oss, då felet ligger i vår förståelseav deras värld, inte i deras förvridna uppfattningar. Även standardexempel på gamla nonsens - debatten om änglar på knappnålshuvuden -vettigt när du inser att teologer inte diskuteradeom fem eller arton skulle passa, men om ett stift kan inrymma enändlig eller ett oändligt antal.
		-- S. J. Gould, "Wide Hats and Narrow Minds"

%
Campus trottoarer finns aldrig som den rakaste linjen mellan två punkter.
		-- M. M. Johnston

%
Jämföra information och kunskap är som att be om fetmaav en gris är mer eller mindre grön än utsedd slagman regeln. "
		-- David Guaspari

%
Kära Freshman,Du vet inte vem jag är och uppriktigt sagt inte bryr sig, menokända för dig vi har något gemensamt. Vi är båda ganskabenägna att misstag. Jag valdes Student Government president frånmisstag, och du kom till skolan här av misstag.
		-- David Guaspari

%
Kära fröken Manners:Min hushållslärare säger att man aldrig får placera sittarmbågarna på bordet. Men jag har läst att en armbåge i mellankurser, är okej. Vilket är korrekt?Gentle läsare:För att besvara undersökningar i ditt hem ekonomiklass, är din lärare korrekt. Fånga på denna princip omutbildning kan vara av ännu större betydelse för dig nu än att lära sigkorrekta aktuella bordsskick, vital som Miss Manners menar att är.
		-- David Guaspari

%
Institutionen ordförande dör aldrig, de bara förlorar sina förmågor.
		-- David Guaspari

%
Visste du University of Iowa stängdes efter någon stal boken?
		-- David Guaspari

%
Inte täppa intellektets slussar med bitar av kunskap om tvivelaktiga användningsområden.
		-- David Guaspari

%
Vet du skillnaden mellan utbildning och erfarenhet? Utbildningär vad du får när du läser det finstilta; erfarenhet är vad du fårnär du inte gör det.
		-- Pete Seeger

%
Tror du att analfabeter få den fulla effekten av alfabetet soppa?
		-- Pete Seeger

%
Utbildning och religion är två saker som inte regleras av tillgång ochefterfrågan. Ju mindre av antingen människor har, desto mindre de vill.
		-- Charlotte Observer, 1897

%
Utbildning är en beundransvärd sak, men det är bra att komma ihåg från tid tilltid att ingenting som är värt att veta kan läras ut.
		-- Oscar Wilde, "The Critic as Artist"

%
Utbildning är att lära sig vad du inte ens vet att du inte vet.
		-- Daniel J. Boorstin

%
Utbildning är en process för gjutning falska pärlor för riktiga svin.
		-- Irwin Edman

%
Utbildning är vad fortlever när vad som har lärt sig har glömts bort.
		-- B. F. Skinner

%
Pedagogiska tv bör absolut förbjudet. Det kan bara ledatill orimligt besvikelse när ditt barn upptäcker att bokstävernai alfabetet inte hoppa upp ur böcker och dansar runt medroyal-blå kycklingar.
		-- Fran Lebowitz, "Social Studies"

%
Vältalighet är logiken i brand.
		-- Fran Lebowitz, "Social Studies"

%
Encyclopedia till salu efter far. Son vet allt.
		-- Fran Lebowitz, "Social Studies"

%
Engineering: "Hur kommer detta arbete?"Science: "Varför kommer detta arbete?"Management: "När kommer detta arbete?"Liberal Arts: "Vill du frites med det?"
		-- Fran Lebowitz, "Social Studies"

%
Även om du inte lära sig tala korrekt engelska, vem ska du taladet till?
		-- Clarence Darrow

%
Överallt jag går jag frågade om jag tror att universitetet kväver författare. Minåsikt är att de inte kväva tillräckligt många av dem. Det finns många en bästsäljaresom kunde ha förhindrats av en bra lärare.
		-- Flannery O'Connor

%
Undersökningar är formidabla även till den bäst förberedda föräven den största idiot kan begära mer den visaste mannen kan svara.
		-- C. C. Colton

%
Erfarenhet är den värsta läraren. Det ger alltid testet först ochinstruktionen efteråt.
		-- C. C. Colton

%
F u cn rd THS u CNT SPL wrth en dm!
		-- C. C. Colton

%
fu cn rd THS, ITN tyg h myxbl cd.
		-- C. C. Colton

%
fu cn rd THS, u cn gt en gd jb n cmptr prgrmmng.
		-- C. C. Colton

%
fu cn rd THS, u r prbbly en LSY spllr.
		-- C. C. Colton

%
Fortune guide till Freshman notetaking:NÄR PROFESSORN SÄGER: Du skriver:Förmodligen den största kvalitet poesi John Milton - född 1608John Milton, som föddes i 1608, är denkombination av skönhet och makt. få harutmärkte honom i användningen av det engelska språket,eller för den delen, i klarhet i versform,"Paradise Lost" sagt att vara den störstaenda dikt som någonsin skrivits. "Aktuella historiker har kommit till de flesta av de problem som nutvivlar hela advantageousness ansiktet USA ärnågra av Roosevelts politik ... direkt spåras tillklumpiga och girighet presidentRoosevelt.... Det är möjligt att vi helt enkelt göra Professor Mitchell är eninte förstå den ryska synvinkel ... kommunist.
		-- C. C. Colton

%
Fjorton år i professor Dodge har lärt mig att man kan argumenteragenialt på uppdrag av någon teori, tillämpas på ett stycke litteratur.Detta är sällan skadlig, eftersom normalt ingen läser dessa essäer.
		-- Robert Parker, quoted in "Murder Ink",  ed. D. Wynn

%
Att gå till kyrkan inte göra en person religiös, inte heller gå i skolangöra en person utbildad, mer än att gå till ett garage gör en person en bil.
		-- Robert Parker, quoted in "Murder Ink",  ed. D. Wynn

%
Bra dag för att undvika polisen. Krypa till skolan.
		-- Robert Parker, quoted in "Murder Ink",  ed. D. Wynn

%
God undervisning är en fjärdedel förberedelse och tre fjärdedelar bra teater.
		-- Gail Godwin

%
Examen liv: Det är inte bara ett jobb. Det är ett AVTAL.
		-- Gail Godwin

%
Doktorander och de flesta professorer är inte smartare än undergrads.De är bara äldre.
		-- Gail Godwin

%
Han som lär sig har en dåre för en mästare.
		-- Benjamin Franklin

%
"Han var en blygsam, godmodig pojke. Det var Oxford som gjorde honom olidlig."
		-- Benjamin Franklin

%
Den som skriver utan felstavade ord har förhindrat en första misstankepå gränserna för sitt stipendium eller, i den sociala världen, hans allmännautbildning och kultur.
		-- Julia Norton McCorkle

%
[Han] tog mig in i hans bibliotek och visade mig sina böcker, som han hadeen komplett uppsättning.
		-- Ring Lardner

%
Högre utbildning hjälper din intjäningsförmåga. Fråga någon college professor.
		-- Ring Lardner

%
Historieböckerna som inte innehåller några lögner är extremt tråkig.
		-- Ring Lardner

%
Historien är ingenting annat än en samling av fabler och onödiga småsaker,belamrad med en massa onödiga siffror och egennamn.
		-- Leo Tolstoy

%
Hur förklarar ni skola till en högre intelligens?
		-- Elliot, "E.T."

%
Jag är en bookaholic. Om du är en anständig person, kommer du inte sälja migen annan bok.
		-- Elliot, "E.T."

%
"Jag är inte säker på vad det är, men en 'F' skulle bara dignify det."
		-- English Professor

%
Jag återkommer detta annars bra att skriva papper till dig eftersom någonhar tryckt rotvälska över det och sätta ditt namn på toppen.
		-- Professor Lowd, English, Ohio University

%
Jag uppskattar det faktum att detta förslag gjordes i all hast, men en del av denmeningar som du skickar ut i världen för att göra ditt arbete för dig ärsölig i krogar eller sover bredvid motorvägen.University of Tennessee på Knoxville
		-- Dr. Dwight Van de Vate, Professor of Philosophy,

%
Jag kom ut från tolv år på college och jag visste inte ens hur man syr.Allt jag kunde göra var konto - Jag kunde inte ens stå för själv.
		-- Firesign Theatre

%
Jag kom till MIT att få en utbildning för mig och ett diplom för min mamma.
		-- Firesign Theatre

%
Jag har gjort detta brev längre än vanligt eftersom jag inte har tid attgöra det kortare.
		-- Blaise Pascal

%
"Jag måste övertyga dig, eller åtminstone snö dig ..."
		-- Prof. Romas Aleliunas, CS 435

%
Jag hörde en definition av en intellektuell, som jag tyckte var mycket intressant:en man som tar fler ord än vad som krävs för att berätta mer än han vet.
		-- Dwight D. Eisenhower

%
Jag respekterar tro, men tvivel är det som ger dig en utbildning.
		-- Wilson Mizner

%
Jag tror att dina åsikter är rimliga, med undantag för den om min mentalainstabilitet.
		-- Psychology Professor, Farifield University

%
"Jag tillbaka denna anmärkning till dig, istället för papper, eftersom det (papperet)närvarande upptar botten av mitt fågelbur. "
		-- English Professor, Providence College

%
Om någon vill bli förödmjukad och beskedet, låt honom bli presidentav Harvard.
		-- Edward Holyoke

%
Om han bara hade lärt sig lite mindre, hur oändligt mycket bättre han kan halärt mycket mer!
		-- Edward Holyoke

%
Om okunnighet är salighet, varför är det inte fler lyckliga människor?
		-- Edward Holyoke

%
Om lite annat, är hjärnan en pedagogisk leksak.
		-- Tom Robbins

%
Om någon hade sagt till mig att jag skulle vara påve en dag, skulle jag ha studerat hårdare.
		-- Pope John Paul I

%
Om högskolor var bättre, om de verkligen hade det, skulle du behöver för att fåpolisen vid grindarna för att hålla ordning i inrushing mångfald. secollege hur vi omintetgöra den naturliga kärlek till lärande genom att lämna den naturligametod för undervisning vad varje önskar att lära sig, och insisterar på att man skalllära sig vad du har ingen smak eller kapacitet för. Högskolan, vilket börvara en plats för härlig arbete, görs motbjudande och ohälsosamma ochunga män lockas till oseriöst nöjen att samla sina jaded sprit.Jag skulle ha studierna valbara. Stipendium ska skapas integenom tvång, utan genom att väcka en ren intresse i kunskap. De visainstruktör åstadkommer detta genom att öppna sina elever justattraktioner studien har för sig själv. Märkningen är ett system för skolor,inte för högskolan; för pojkar, inte för män; och det är en ungracious arbete attsätta på en professor.
		-- Ralph Waldo Emerson

%
Om sanningen är skönhet, hur kommer ingen har sitt hår gjort i biblioteket?
		-- Lily Tomlin

%
Om vi ​​talade ett annat språk, skulle vi uppfattar en något annorlunda värld.
		-- Wittgenstein

%
Om medan du är i skolan, det finns en brist på kvalificerad personalinom ett visst område, så med den tid du examen med nödvändigkvalifikationer, är det fältets arbetsmarknaden glutted.
		-- Marguerite Emmons

%
Om du är för upptagen för att läsa, då du är för upptagen.
		-- Marguerite Emmons

%
Om du inte kan läsa detta, skyller en lärare.
		-- Marguerite Emmons

%
Om du motstå läsa vad du inte håller med, hur kommer du någonsin fådjupare insikter i vad du tror? De saker mest läsvärdär just de som utmanar våra övertygelser.
		-- Marguerite Emmons

%
Om du tror att utbildning är dyrt, prova okunnighet.
		-- Derek Bok, president of Harvard

%
Om du tog alla elever som kände sover i klassen och lade dem slut påDärför skulle de vara mycket mer bekväm.
		-- "Graffiti in the Big Ten"

%
"Om du förstår vad du gör, du är inte lära sig något."
		-- A. L.

%
Okunnighet är aldrig omodernt. Det var på modet i går, är detrasa idag, och det kommer att ange takten i morgon.
		-- Franklin K. Dane

%
Okunnighet är när man inte vet någonting och någon hittar den ut.
		-- Franklin K. Dane

%
Okunnighet måste verkligen vara salighet eller skulle det inte finnas så många människorså beslutsamt fullfölja den.
		-- Franklin K. Dane

%
Analfabet? Skriv idag, gratis hjälp!
		-- Franklin K. Dane

%
I en skog en räv stöter en liten kanin, och säger: "Hej,Junior, vad håller du på med? ""Jag skriver en avhandling om hur kaniner äter rävar", sadekanin."Kom nu, kompis kanin, du vet att det är omöjligt! Ingenpublicerar sådant skräp! ""Nå, följ mig och jag ska visa dig."De båda går in i kaninens bostad och efter en stundkanin framträder med en nöjd uttryck i ansiktet. Kommer tillsammans envarg. "Hej, lilla kompis, vad gör vi dessa dagar?""Jag skriver 2'nd kapitlet i min avhandling om hur kaniner slukarvargar. ""Är du galen? Var är din akademisk hederlighet?""Kom med mig och jag ska visa dig."Liksom tidigare kommer kaninen ut med en nöjd blick på hans ansikteoch en examen i sin tass. Slutligen, kameran panorerar i kaninen grottaoch, som alla skulle ha gissat vid det här laget, ser vi en genomsnittlig utseende, storlejon, sittande, plocka sina tänder och rapningar, bredvid några furry, blodigresterna av varg och räv.Sensmoralen: Det är inte innehållet i avhandlingen som ärviktigt - det är din PhD rådgivare som verkligen räknas.
		-- Franklin K. Dane

%
I Kalifornien, Bill Honig, vicevärden av offentlig anvisning, sade hantrodde allmänheten bör ha en röst i att definiera vad en utmärktlärare bör veta. "Jag skulle inte lämna definitionen av matematik," Dr Honigsa, "upp till matematiker."
		-- The New York Times, October 22, 1985

%
I stället för att ge pengar till hittade högskolor för att främja lärande, varför intede passerar en konstitutionstillägg som förbjuder någon från lärandenågot? Om det fungerar lika bra som förbud mot en gjorde, varför i femår skulle vi ha smartaste ras av människor på jorden.
		-- The Best of Will Rogers

%
Iowa State - gymnasiet efter gymnasiet!
		-- Crow T. Robot

%
Det har sagts [av Anatole France], "det är inte genom att roa sigatt man lär sig ", och som svar:" det är * ____ bara * av roar sig attman kan lära sig. "
		-- Edward Kasner and James R. Newman

%
Det har länge varit ett föremål för vår folklore att för mycket kunskap eller skicklighet,eller särskilt fulländad kompetens, är en dålig sak. Det avhumaniserar dem somuppnå det, och gör det svårt deras handel med bara vanlig folk, i vilkagamla goda sunt förnuft inte har utplånats av ren bok lärande eller fantasiföreställningar. Denna populära villfarelse blomstrar nu mer än någonsin, för vi är allainfekterade med det i skolan, där pedagoger har förhöjda det frånfolklore artikel av Tro. Det ökar deras självkänsla och ljusarederas arbete genom att tillhandahålla teoretisk motivering för att besluta attuppskattning, eller även enkla medvetenhet, är mer att uppskattad än kunskap,och rör (till sig själv och andra), mer än skicklighet, där minimikompetens kommer att vara helt tillräckligt.
		-- The Underground Grammarian

%
Det är en djupt felaktig truism, upprepas av alla kopierings-böcker ochav framstående personer när de gör tal, att vi bör odlaför vana att tänka på vad vi gör. Den exakta motsatsen ärfall. Civilization framsteg genom att förlänga antalet viktiga operationersom vi kan utföra utan att tänka på dem. Verksamheten tanke ärsom kavalleri avgifter i strid - de är strängt begränsade i antal, dekräver nya hästar och får endast ske till avgörande ögonblick.
		-- Alfred North Whitehead

%
Det är grad examen tid ...DATAVETENSKAPInuti skrivbordet hittar du en lista över DEC / VMS operativsystemsystemet i IBM 1710 maskinkod. Visa vilka förändringar som krävs för att omvandladenna kod i en UNIX Berkeley 7 operativsystem. Bevisa att dessa korrigeringar ärbuggfri och fungera korrekt. Du bör få minst 150% effektivitet inya systemet. (Du bör inte ta mer än 10 minuter på denna fråga.)MATEMATIKOm X är lika med PI gånger R ^ 2, konstruera en formel som visar hur lång tiddet skulle ta en brand myra att borra ett hål genom en dill pickle, omlängd omkrets förhållandet mellan myran till pickle var 98,17: 1.ALLMÄNBILDNINGBeskriv universum. Ge tre exempel.
		-- Alfred North Whitehead

%
Det är grad examen tid ...MEDICINDu har försetts med ett rakblad, en bit gasbinda, och enflaska Scotch. Ta bort blindtarmen. Suturera inte förrän ditt arbete harinspekterats. (Du har 15 minuter.)HISTORIABeskriv historia påvedömet från sitt ursprung till idagdag, framför allt vad, men inte uteslutande, på dess sociala, politiska,ekonomiska, religiösa och filosofisk påverkan på Europa, Asien, Amerika, ochAfrika. Vara korta, koncisa och specifik.BIOLOGISkapa liv. Uppskatta skillnaderna i efterföljande mänsklig kulturom denna form av liv hade skapats 500 miljoner år sedan eller tidigare, medsärskild uppmärksamhet åt dess troliga inverkan på engelska parlamentariska systemet.
		-- Alfred North Whitehead

%
Det är inte, det är inte är inte, och det är det, inte dess, om du menar detär. Om du inte gör det, är det dess. Även då det är hennes. Det är inte hennes talet. Detär inte vår är antingen. Det är vår, och likaså din och deras.
		-- Oxford University Press, Edpress News

%
Joe Cool tillbringar alltid de två första veckorna på college segling sin frisbee.
		-- Snoopy

%
Lärda män är cisterner kunskap, inte fountainheads.
		-- Snoopy

%
Att lära på vissa skolor är som att dricka ur en brandslang.
		-- Snoopy

%
Att lära utan tanke är arbete förlorad;tanken utan lärande är farlig.
		-- Confucius

%
Kanske är inte inte så korrekt, men jag märker att massor av folk som inte äranvänder inte inte Eatin väl.
		-- Will Rogers

%
De flesta seminarierna har ett lyckligt slut. Alla är glada när de är över.
		-- Will Rogers

%
Min far, en god man, berättade, "förlorar aldrig din okunnighet, du kan inteErsätt den."
		-- Erich Maria Remarque

%
Aldrig har så många förstått så lite om så mycket.
		-- James Burke

%
Låt aldrig din skolgång störa din utbildning.
		-- James Burke

%
Ingen disciplin någonsin fordrar att tvinga närvaro på föreläsningar som ärverkligen värt att delta.
		-- Adam Smith, "The Wealth of Nations"

%
Oavsett vem du är, kan en del forskare visa den stora idé du hadevar hade någon före dig.
		-- Adam Smith, "The Wealth of Nations"

%
Inte konstigt att du är trött! Du förstod så mycket idag.
		-- Adam Smith, "The Wealth of Nations"

%
Normalt våra regler är stela; vi tenderar att diskretion, om av någon annan anledningän självförsvar. Vi rekommenderar aldrig någon av våra studenter, även om viglatt ge information till dem som har misslyckats sina kurser.
		-- Jack Vance, "Freitzke's Turn"

%
Inte bara är detta obegripligt, men bläcket är ful och papperär från fel typ av träd.Jag ser fram emot att arbeta med dig på detta nästa år.
		-- Professor, Harvard, on a  senior thesis.

%
`O 'NIVÅ motkulturTimewarp tillåtet: 3 timmar. Inte scrawl situationalist graffiti imarginaler eller stub dina samlade i inkwells. Orange kan bäras. Krediterakommer att ges till kandidater som själv aktualisera.(1) Jämför och kontrast Pink Floyd med Black Sabbath och säga varförvarken har gatan trovärdighet.(2) "Även Buddha skulle ha varit svårt att nå Nirvana hukpå en ångvält väg. "Tänk på dialektik inre sanningoch innerstaden.(3) Diskutera grad av besvär som deltar i paranoia om att sugasin i ett svart hål.(4) "The egomaniac s Liberation Front var ett gäng revisionistripoff handlare. "Kommentera denna förolämpning.(5) står för bristen på hänvisningar till brunt ris i Dylans texter.(6) "Castenada var lite av en bozo." Hur långt är detta en rättvis summeringav västra dualism?(7) Hermann Hesse var en Fiskarna. Diskutera.
		-- Professor, Harvard, on a  senior thesis.

%
"OK, nu ska vi titta på fyra dimensioner på tavlan."
		-- Dr. Joy

%
OK, så du är en Ph.D. Bara inte röra någonting.
		-- Dr. Joy

%
Man kan inte göra en omelett utan att knäcka ägg - men det är fantastiskthur många ägg man kan bryta utan att göra en anständig omelett.
		-- Professor Charles P. Issawi

%
PERIFRAS är att sätta saker i en rondell sätt. "Kostnaden kan varauppemot en siffra snarare under 10m #. "är en PERIFRAS för Kostnaden kan varanästan 10m #. "I Paris finns regerar en total avsaknad av riktigt pålitligtnyheter "är en PERIFRAS för Det finns ingen tillförlitlig nyheter i Paris." Sällan gör"Lilla Summer dröja fram till november, men ibland sin vistelse har varitförlängdes till ganska sent i årets näst sista månaden "innehåller enPERIFRAS för november, och en annan för dröjer. "Svaret är inegativ "är en PERIFRAS för Nej" Gjordes mottagaren av "är enPERIFRAS för Presenterades med. Den PERIFRAS stil är knappast möjligtpå någon större skala utan mycket användning av abstrakta substantiv som "bas,fall tecken, Connexion, brist, beskrivning, varaktighet, ram, brist,natur, referens, avseende respekt ". Förekomsten av abstrakta substantiv är enbevis på att abstrakt tänkande har skett; abstrakt tänkande är ett tecken påciviliserade människan; och det har kommit om att PERIFRAS och civilisationav många anses vara oskiljaktiga. Dessa goda människor känner att det finns ett nästanoanständigt nakenhet, en återgång till barbari, att säga Inga nyheter är goda nyheteri stället för "Frånvaron av intelligens är en indikation på tillfredsställandeutvecklingen. "
		-- Fowler's English Usage

%
"Plaese porrf Raed."
		-- Prof. Michael O'Longhlin, S.U.N.Y. Purchase

%
Praxis är den bästa av alla lärare.
		-- Publilius

%
Princeton smak är söt som en jordgubbstårta. Harvards är en subtilsmak, som whisky, kaffe, eller tobak. Det kan även vara en dålig vana, förallt jag vet.
		-- Prof. J. H. Finley '25

%
Professor Gorden Newell kastade en annan shutout i förra veckans Chem Eng. 130halva tiden. Än en gång en elev inte fått en enda punkt på sin examen.Newell har nu kastade 5 shutouts detta kvartal. Newells tjänade tenta genomsnittligahar nu sjunkit till en fenomenal 30%.
		-- Prof. J. H. Finley '25

%
Läsning tänker med någon annans huvud i stället för en egen.
		-- Prof. J. H. Finley '25

%
Läsning är att sinnet vad motion är för kroppen.
		-- Prof. J. H. Finley '25

%
Reporter: "Hur kunde du skolan när du växte upp, Yogi?"Yogi Berra: "Closed."
		-- Prof. J. H. Finley '25

%
Regler för god Grammar # 4.(1) Använd inte några dubbla negativ.(2) Gör varje pronomen överens med sina föregångare.(3) Gå klausuler bra, som en förening ska.(4) Om dem meningen fragment.(5) När dinglande, titta på dina participles.(6) Verb har fått att komma överens med sina undersåtar.(7) Bara mellan dig och jag är viktigt fall.(8) Skriv inte köras på straff när de är svåra att läsa.(9) Använd inte kommatecken, som inte är nödvändiga.(10) Försök att aldrig dela infinitiv.(11) Det är viktigt att använda apostrof är korrekt.(12) Korrekturläs ditt skrivande att se om du några ord ur.(13) Korrekt speling är viktigt.(14) En preposition är något du aldrig avsluta en mening med.(15) Även om en transcen ordförråd är lovvärd, måste man vara för evigtförsiktig så att den beräknade målet för kommunikation intebli ensconsed i dunkel. Med andra ord, undfly förvirring.
		-- Prof. J. H. Finley '25

%
Smartness körs i min familj. När jag gick i skolan var jag så smart minlärare var i min klass i fem år.
		-- George Burns

%
Vissa forskare är som åsnor, de bara bära en massa böcker.
		-- Folk saying

%
"Speed ​​är subsittute fo noggrannhet."
		-- Folk saying

%
Stavning är en lossed konst.
		-- Folk saying

%
Plötsligt inser professor Liebowitz han har kommit till seminarietutan hans anka ...
		-- Folk saying

%
Lärarna har klass.
		-- Folk saying

%
"A" är för innehåll, är "minus" för att inte skriva det. Inte någonsin göradetta i mina ögon igen.
		-- Professor Ronald Brady, Philosophy, Ramapo State College

%
Väckarklockan som är högre än Guds egen tillhör rumskamrat medden tidigaste klassen.
		-- Professor Ronald Brady, Philosophy, Ramapo State College

%
Den genomsnittliga Ph.D avhandling är ingenting annat än överföring av ben frånen graveyard till en annan.
		-- J. Frank Dobie, "A Texan in England"

%
Den avocation att bedöma misslyckanden bättre män kan vridasi en bekväm försörjning, förutsatt att du backa upp det med en Ph.D.
		-- Nelson Algren, "Writers at Work"

%
"Det bästa för att vara ledsen", svarade Merlin, börjar puffoch slag, "är att lära sig något. Det är det enda som aldrig misslyckas.Du kan åldras och darrande i dina anatomies, kan du ligga vaken pånatt lyssnar på sjukdom i dina ådror, kan du missar din enda kärlek,du kan se världen om du drabbats av onda galningar, eller kännaära trampade i kloakerna av baser sinnen. Det finns bara en sak fördet då - att lära sig. Läs om varför världen viftar och vad viftar det. Det ärdet enda som sinnet aldrig kan uttömma aldrig stöta aldrig varatorterad av, aldrig rädd eller misstro, och aldrig drömma om att beklaga. Inlärningär det enda för dig. Titta vad en hel del saker som finns att lära. "
		-- T. H. White, "The Once and Future King"

%
Hjärnan är en underbar organ; det börjar arbeta så fort du får upppå morgonen, och inte sluta förrän du kommer till skolan.
		-- T. H. White, "The Once and Future King"

%
College examen presenteras med en fårskinn för att täcka hansintellektuell nakenhet.
		-- Robert M. Hutchins

%
Slutet av världen kommer att ske vid 03:00, på fredag, medsymposium att följa.
		-- Robert M. Hutchins

%
Framtiden är en tävling mellan utbildning och katastrof.
		-- H. G. Wells

%
Det viktiga är inte att stoppa förhör.
		-- H. G. Wells

%
Mannen som aldrig har piskade aldrig har lärt.
		-- Menander

%
Det enda som erfarenheten lär oss är att erfarenheten lär oss ingenting.
		-- Andre Maurois (Emile Herzog)

%
Det enda vi lär av historien är att vi inte lär.Att män inte lär mycket av historien är det viktigaste av alltde lärdomar som historien har att lära.Vi lär oss av historien som vi inte lär av historien.HISTORIA: Papa Hegel han säger att allt vi lär av historien är att vi läringenting av historien. Jag känner folk som inte ens kan lära av vad som händeden här morgonen. Hegel måste ha tagit ett längre perspektiv.
		-- Chad C. Mulligan, "The Hipcrime Vocab"

%
Det enda vi lär av historien är att vi lär oss ingenting av historien.Jag vet killar kan inte lära från igår ... Hegel måste ta ett längre perspektiv.
		-- John Brunner, "Stand on Zanzibar"

%
Problemet med doktorander, i allmänhet, är att de haratt sova med några dagars mellanrum.
		-- John Brunner, "Stand on Zanzibar"

%
Förhållandet av läs- och skrivkunnighet för att analfabetism är en konstant, men numera denanalfabeter kan läsa.
		-- Alberto Moravia

%
Det verkliga syftet med böcker är att fånga sinnet till att göra sitt eget tänkande.
		-- Christopher Morley

%
"Studenten i fråga utför minimalt för hans jämnåriga ochär en framväxande underachiever. "
		-- Christopher Morley

%
Summan av intelligens världen är konstant. Befolkningen är,naturligtvis, växer.
		-- Christopher Morley

%
De sunlights skiljer sig åt, men det finns bara ett mörker.
		-- Ursula K. LeGuin, "The Dispossessed"

%
Testet av en förstklassig intelligens är förmågan att hålla två motsattaidéer i sinnet samtidigt och ändå behålla förmågan att fungera.
		-- F. Scott Fitzgerald

%
De tre bästa sakerna med att gå i skolan är juni, juli och augusti.
		-- F. Scott Fitzgerald

%
The Tree of Learning bär den ädlaste frukt, men ädel frukt smakar illa.
		-- F. Scott Fitzgerald

%
USA är så enorm, och så många är dess skolor, högskolor och religiösaseminarier, många ägnas åt särskilda religiösa övertygelse som sträcker sig frånoortodoxa till dotty, att vi knappast kan undra på sin vilket ger en merbounteous skörd av gobbledegook än resten av världen tillsammans.
		-- Sir Peter Medawar

%
Världen kommer till ett slut! Omvänd er och återlämna dessa biblioteksböcker!
		-- Sir Peter Medawar

%
Världen är full av människor som aldrig har, sedan barndomen, träffade enöppna dörren med ett öppet sinne.
		-- E. B. White

%
Det finns inga svar, bara korsreferenser.
		-- Weiner

%
Detta är den typ av engelska med som jag inte kommer att sätta.
		-- Winston Churchill

%
De som utbildar barn väl är mer att hedras än föräldrarna, fördessa bara gav liv, de konsten att leva väl.
		-- Aristotle

%
Tid är en stor lärare, men tyvärr det dödar alla sina elever.
		-- Hector Berlioz

%
Att anklaga andra för sina egna olyckor är ett tecken på brist på utbildning.Att anklaga sig själv visar att en utbildning har påbörjats. Anklaga varkensjälv eller andra visar att en utbildning är klar.
		-- Epictetus

%
Att craunch en silkesapa.
		-- Pedro Carolino, "English as She is Spoke"

%
Att undervisa är att lära sig två gånger.
		-- Joseph Joubert

%
Att undervisa är att lära sig.
		-- Joseph Joubert

%
Försök att inte ha en god tid ... Detta är tänkt att vara lärorikt.
		-- Charles Schulz

%
Att försöka få en utbildning här är som att försöka få en drink från en brandslang.
		-- Charles Schulz

%
Universiteten är platser för kunskap. Den förstaårselev varje få litein med dem, och de äldre tar ingen bort, så kunskap ackumuleras.
		-- Charles Schulz

%
Universitets politik är ond just eftersom insatserna är så små.
		-- C. P. Snow

%
Walt: Pappa, vad är gradvis skolan?Garp: Gradvis skolan?Walt: Ja. Mamma säger att hennes arbete är roligare nu när hon undervisargradvis skola.Garp: Oh. Tja, är gradvis skola någonstans du gå och gradvista reda på att du inte vill gå till skolan längre.
		-- The World According To Garp

%
"Vi kräver fast definierade områden av tvivel och osäkerhet!"
		-- Vroomfondel

%
Vi vet nästan ingenting om nästan allt. Det är inte nödvändigtatt veta varifrån universum; Det är nödvändigt att vill veta.Civilisation beror inte på någon särskild kunskap, men om dispositionerlängta kunskap.
		-- George Will

%
Vi är fantastiskt otroligt synd om alla dessa extremt orimligtsaker som vi gjorde. Jag kan bara göra gällande att min enkla, knappt kännande vänoch jag är underprivilegierade, berövade och även studenter.
		-- Waldo D. R. Dobbs

%
"Vi kör ut adjektiv för att beskriva vår situation. Vihade kris, sedan gick vi in ​​i kaos, och nu vad vi kallar detta gör "sa?Nicaraguas ekonomen Francisco Mayorga, som har en doktorsexamen från Yale.New Yorker kommentar:Vid Harvard skulle de kallar det ett substantiv.
		-- The Washington Post, February, 1988

%
Vad gör utbildning ofta gör? Det gör ett rakt snitt dike av enfri slingrande bäck.
		-- Henry David Thoreau

%
Vad jag gjorde under min höstterminenPå den första dagen av min hösttermin, jag fick upp.Sedan gick jag till biblioteket för att hitta ett uppsatsämne.Sen hängde framför Dover.På den andra dagen av min hösttermin, jag fick upp.Sedan gick jag till biblioteket för att hitta ett uppsatsämne.Sen hängde framför Dover.På den tredje dagen av min hösttermin, jag fick upp.Sedan gick jag till biblioteket för att hitta ett uppsatsämne.Jag hittade en avhandling ämne:Hur att hålla folk från att hänga ut framför Dover.
		-- Sister Mary Elephant, "Student Statement for Black Friday"

%
Varför tror du att forskarskolan är tänkt att tillfredsställa?
		-- Erica Jong, "Fear of Flying"

%
Vad passerar för optimism är oftast effekten av en intellektuell fel.
		-- Raymond Aron, "The Opium of the Intellectuals"

%
Vad vi inte förstår att vi inte har.
		-- Goethe

%
Vad är sidan en, ett förebyggande anfall?
		-- Professor Freund, Communication, Ramapo State College

%
När jag var i skolan, jag var otrogen mot min metafysik examen: Jag tittade insjäl pojke som sitter bredvid mig.
		-- Woody Allen

%
När någon säger, "teoretiskt" de egentligen "inte riktigt."
		-- Dave Parnas

%
Var kan jag hitta tid för att inte läsa så många böcker?
		-- Karl Kraus

%
"Vem är du?" sade han, för han hade varit på kvällskurs.
		-- George Ade

%
Skulle inte meningen "Jag vill sätta ett bindestreck mellan orden fiskoch och och och och Chips i min fisk-och-chips tecken "har varit tydligare omcitattecken hade placerats före fisk och mellan fisk och och ochoch och och och och och och och och och och och och och och och och ochChips, liksom efter Chips?
		-- George Ade

%
Du kan inte förvänta sig en pojke att vara ond tills han har varit en bra skola.
		-- H. H. Munro

%
Du behöver inte tänka för hårt när du pratar med lärare.
		-- J. D. Salinger

%
Du kanske har hört att en dekanus är att lärare som brandpost är en hund.
		-- Alfred Kahn

%
"Du bör utan tvekan, pund din skrivmaskin i en plowshare,dina papper till gödsel och ange jordbruk "
		-- Business Professor, University of Georgia

%
Din utbildning börjar där det som kallas din utbildning är över.
		-- Business Professor, University of Georgia

%
