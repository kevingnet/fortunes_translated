VägenDet sätt som kan upplevas är inte sant;Den värld som kan konstrueras är inte verkligt.Vägen visar allt som händer och kan hända;Världen representerar allt som existerar och kan förekomma.Att uppleva utan abstraktion är att känna världen;Att uppleva med abstraktion är att känna världen.Dessa två upplevelser är oskiljbara;Deras konstruktion skiljer sig men deras effekt är densamma.Bortom grinden erfarenhet flyter Way,Som är allt större och mer subtila än världen.
		-- Lao Tse, "Tao Te Ching"

%
AbstraktionNär skönhet abstraheradeDå fulhet har antytts;När bra abstraherasSedan det onda har antytts.Så levande och döda sammandrag från naturen,Svårt och lätt abstraherade från framsteg,Långa och korta sammandrag från kontrast,Högt och lågt abstraherade från djupet,Sång och tal sammandrag från melodi,Efter och före abstraherade från sekvens.Den vise erfarenheter utan abstraktion,Och åstadkommer utan åtgärd;Han accepterar ebb och flod av saker,Vårdar dem, men inte äger dem,Och lever, men inte bo.
		-- Lao Tse, "Tao Te Ching"

%
utan åtgärdInte berömma värdig förhindrar påstående,Inte esteeming värdefulla förhindrar stöld,Inte visa vackra förhindrar önskan.På detta sätt den vise styr folk:Tömma sina sinnen,Fylla sina magar,Försvagar deras ambitioner,Och stärka deras ben.Om människor saknar kunskap och lustDå de inte kan agera;Om inga åtgärder vidtasHarmoni återstår.
		-- Lao Tse, "Tao Te Ching"

%
GränslösVägen är en gränslös kärl;Används av sig själv, är det inte fylls av världen;Det kan inte skäras, knutna, nedtonade eller stillad;Dess djup är dolda, allestädes närvarande och evigt;Jag vet inte varifrån det kommer,Det kommer före naturen.
		-- Lao Tse, "Tao Te Ching"

%
NaturNaturen är inte snäll,Den behandlar allt opartiskt.Sage är inte snäll,Och behandlar alla människor opartiskt.Naturen är som en bälg,Tom, men aldrig upphör sin försörjning.Ju mer den rör sig, ger desto mer;Så den vise bygger på erfarenhetOch kan inte vara uttömda.
		-- Lao Tse, "Tao Te Ching"

%
ErfarenhetErfarenhet är en flodbädd,Dess källa dold, alltid flyter:Dess entré, roten av världen,Vägen rör sig inom det:Utnyttja det; det kommer inte att köras torr.
		-- Lao Tse, "Tao Te Ching"

%
KomplettNaturen är fullständig eftersom det inte tjänar själv.Den vise placerar sig själv efter och finner sig inför,Ignorerar hans önskan och befinner sig innehåll.Han är komplett eftersom han inte tjänar själv.
		-- Lao Tse, "Tao Te Ching"

%
VattenDet bästa av människan är som vatten,Vilket gynnar alla ting, och inte brottas med dem,Som flyter på platser som andra förakt,Om det är i harmoni med vägen.Så vis:Bor inom natur,Tänker inom den djupa,Ger inom opartiskhet,Talar inom tillit,Reglerar inom ordning,Hantverk inom förmåga,Agerar inom tillfälle.Han har inte påstått, och ingen hävdar mot honom.
		-- Lao Tse, "Tao Te Ching"

%
Gå i pensionFyll en kopp till dess brädden och det är lätt spills;Mildra ett svärd till dess svåraste och det är lätt bryts;Samla den största skatten och det är lätt stulen;Anspråk på kredit och ära och du enkelt falla;Dra dig tillbaka när ditt syfte uppnås - detta är naturligt.
		-- Lao Tse, "Tao Te Ching"

%
HarmoniOmfamna vägen, blir du anammat;Andas försiktigt, blir du nyfödda;Rensa ditt sinne, du blir klar;Vårda dina barn, du blir opartisk;Öppna ditt hjärta, du blir accepterad;Acceptera världen, omfamna dig vägen.Bäring och vårda,Skapa men inte äga,Ge utan att kräva,Detta är harmoni.
		-- Lao Tse, "Tao Te Ching"

%
verktygTrettio ekrar möts vid en skeppet;På grund av hålet vi kan använda hjulet.Lera formas till ett kärl;På grund av den ihåliga vi får använda koppen.Väggar är uppbyggda kring en härd;På grund av dörrarna kan vi använda huset.Således verktyg kommer från vad som finns,Men använda från vad som inte fungerar.
		-- Lao Tse, "Tao Te Ching"

%
ÄmneFör mycket färg förblindar ögat,För mycket musik deafens örat,För mycket smak dämpar gommen,För stort spel Maddens sinnet,För mycket önskan tårar hjärtat.På detta sätt den vise bryr sig om människor:Han ger magen, inte för alla sinnen;Han ignorerar abstraktion och håller fast vid ämnet.
		-- Lao Tse, "Tao Te Ching"

%
SjälvBåde ris och ros orsaka oro,För de föra människor hopp och fruktan.Syftet med hopp och fruktan är själv -Ty utan själv, vem kan lycka och katastrof inträffar?Därför,Vem som skiljer sig från världen kan ges i världen,Men som betraktar sig själv som världens kan acceptera världen.
		-- Lao Tse, "Tao Te Ching"

%
MysteriumTittat på men kan inte ses - är den under form;Lyssnade på men kan inte höras - det är under ljud;Hölls men kan inte röras - är den under känsla;Dessa depthless saker undgå definition,Och blanda i ett enda mysterium.I sin stigande det finns inget ljus,I sin faller det finns inget mörker,En kontinuerlig tråd bortom beskrivning,Foder vad som inte finns;Dess form formlös,Dess bild ingenting,namn tystnad dess;Följ den, det har ingen back,Möta det, har den ingen ansikte.Delta i närvarande för att ta itu med det förflutna;Således du förstå kontinuiteten på vägen,Som är dess väsen.
		-- Lao Tse, "Tao Te Ching"

%
UpplysningDen upplysta besitter förståelseSå djup att de inte kan förstås.Eftersom de kan inte förståsJag kan bara beskriva deras utseende:Försiktig som en korsning tunn is,Inte bestämt som en omgiven av fara,Modest som en som är en gäst,Gränslös som smältande is,Äkta som unshaped trä,Bred som en dal,Smidig som grumligt vatten.Vem stillar vattnet att leran får avgöra,Som försöker sluta att han kan resa vidare,Som önskar mindre än vad som kan sippra ut,Sönderfaller, men kommer inte att förnya.
		-- Lao Tse, "Tao Te Ching"

%
Förfall och förnyelseTöm själv helt;Omfamna perfekt fred.Världen kommer att stiga och flytta;Se den återgå till vila.Alla blomstrande sakerKommer tillbaka till sin källa.Denna avkastning är fredlig;Det är flödet av naturen,Ett evigt förfall och förnyelse.Acceptera detta ger upplysning,Att ignorera detta medför elände.Som accepterar naturens flöde blir all-cherishing;Att all-cherishing han blir opartisk;Att vara opartisk han blir storsint;Att vara storsint han blir naturligt;Att vara naturligt att han blir ett med vägen;Att vara ett med hur han blir odödlig:Även om hans kropp kommer att förfalla, vägen kommer inte.
		-- Lao Tse, "Tao Te Ching"

%
linjalerDe bästa härskare är knappast kända av sina undersåtar;Det näst bästa är älskade och prisade;Nästa befaras;Nästa föraktade:De har ingen tro på deras folk,Och deras folk blir otrogen dem.När de bästa härskare uppnår sitt syfteSina undersåtar göra anspråk på prestation som sin egen.
		-- Lao Tse, "Tao Te Ching"

%
HyckleriNär vägen glömsTull och rättvisa visas;Då kunskap och visdom födsTillsammans med hyckleri.När harmoniska relationer upplösaDå respekt och hängivenhet uppstår;När en nation faller till kaosDå lojalitet och patriotism föds.
		-- Lao Tse, "Tao Te Ching"

%
FörenklaOm vi ​​kunde kassera kunskap och visdomDå folk skulle dra hundrafalt;Om vi ​​kunde kasta plikt och rättvisaDå skulle harmoniska relationer bildas;Om vi ​​kunde kasta knep och vinstDå avfall och stöld skulle försvinna.Men sådana åtgärder behandla bara symptomOch så de är otillräckliga.Människor behöver personliga åtgärder:Avslöja din nakna själv och omfamna din ursprungliga natur;Binda egenintresse och styra din ambition;Glöm dina vanor och förenkla dina affärer.
		-- Lao Tse, "Tao Te Ching"

%
VandrandeVad är skillnaden mellan samtycke och förnekande?Vad är skillnaden mellan vackra och fula?Vad är skillnaden mellan skräckinjagande och rädd?Folk är glada, som om på en magnifik festEller leker i parken vid våren,Men jag är lugn och vandra,Som en nyfödd innan den lär sig att le,Ensam, utan sanna hem.Folket har i överflöd,Där jag har ingenting,Och mitt hjärta är dumt,Rörig och grumlig.Människorna är ljusa och säker,Där jag är svag och förvirrad;Människorna är smarta och kloka,Där jag är tråkig och okunniga;Mållöst som en våg drivande över havet,Bifogat till ingenting.Folk är upptagen med syfte,Där jag är opraktiskt och grov;Jag delar inte folkens bekymmerMen jag är trött på naturens bröst.
		-- Lao Tse, "Tao Te Ching"

%
AccepteraHarmoni är bara att följa vägen.Vägen är utan form eller kvalitet,Men uttrycker alla former och kvaliteter;Vägen är dold och blandar,Men uttrycker hela naturen;Vägen är oföränderliga,Men uttrycker all rörelse.Beneath sensation och minneVägen är källan till hela världen.Hur kan jag förstå källan av världen?Genom att acceptera.
		-- Lao Tse, "Tao Te Ching"

%
HemAcceptera och du blir hela,Bend och du räta,Töm och du fyller,Förfall och du förnyar,Vill och du förvärva,Uppfylla och du blir förvirrad.Den vise accepterar världenSom världens accepterar vägen;Han visar inte sig själv, så syns tydligt,Inte rättfärdiga sig själv, så är erkänd,Skryter inte, så krediterasInte stolthet själv, så uthärdar,Har inte påstått, så ingen kämpa mot honom.Den gamle sade, "Acceptera och du blir helt",När hela, är världen som ditt hem.
		-- Lao Tse, "Tao Te Ching"

%
OrdNaturen säger endast ett fåtal ord:Hög vinden inte länge,Inte heller kraftiga regn.Om naturens ord inte vararVarför skulle de av människan?Som accepterar harmoni blir harmonisk.Som accepterar förlust, förloras.För som accepterar harmoni, harmonierar med honom på vägen,Och som accepterar förlust, kan vägen inte hitta.
		-- Lao Tse, "Tao Te Ching"

%
FlathetRäta själv och du kommer inte stå stadigt;Visa dig själv och du kommer inte att tydligt;Motivera dig själv och du kommer inte att respekteras;Marknadsföra dig själv och du kommer inte bli trodd,Stolthet själv och du kommer inte att uthärda.Dessa beteenden är slösaktig, överseende,Och så de locka onåd;Harmoni undviker dem.
		-- Lao Tse, "Tao Te Ching"

%
Beneath abstraktionDet är ett mysterium,Under abstraktion,Tyst, depthless,Ensam, oföränderlig,Ubiquitous och vätska,Moder natur.Den har inget namn, men jag kallar det "vägen";Det har ingen gräns, men jag kallar det "gränslösa".Att vara obegränsad, flyter bort för alltid;Flödande bort för evigt, återgår den till mig själv:Vägen är gränslös,Så naturen är gränslös,Så världen är obegränsade,Och så är jag gränslös.För jag abstraherade från världen,Världen från naturen,Natur från vägen,Och vägen från vad som är under abstraktion.
		-- Lao Tse, "Tao Te Ching"

%
LugnaGravity är källan av lätthet,Lugn, befälhavare brådska.En ensamstående resenär kommer resa hela dagen, vakar över sintillhörigheter;Enda säkra i sin egen säng kan han förlora dem i sömnen.Så kaptenen på en stor fartyg bör inte agera lätt eller hastigt.Agera lätt, förlorar han syn på världen,Agera hastigt, förlorar han kontrollen över sig själv.Kaptenen kan inte behandla hans stora fartyg som en liten båt;Snarare än glitter som jadeHan måste stå som sten.
		-- Lao Tse, "Tao Te Ching"

%
FulländningDen perfekta resenären lämnar inget spår som skall följas;Den perfekta högtalaren lämnar ingen fråga som måste besvaras;Den perfekta revisor lämnar ingen fungerande slutföras;Den perfekta behållare lämnar inga lås att stängas;Den perfekta knut lämnar inget slut att ravelled.Så salvia vårdar alla mänOch överger ingen.Han accepterar alltOch avvisar ingenting.Han deltar i minsta detalj.För den starka måste styra svaga;Den svaga är råvara till de starka.Om guiden inte respekteras,Eller materialet inte vårdas,Förvirring kommer att resultera, oavsett hur duktig man är.Detta är hemligheten bakom perfektion:När obehandlat trä är huggen, blir det ett verktyg;När en man är anställd, blir han ett verktyg;Den perfekta snickare lämnar ingen ved att lyftas.
		-- Lao Tse, "Tao Te Ching"

%
PassandeMed hjälp av manliga, vara kvinna,Att vara ingången till världen,Du omfamna harmoniOch bli som en nyfödd.Med hjälp av styrka, att vara svag,Är roten av världen,Du fullständig harmoniOch bli lika unshaped trä.Med hjälp av ljus, som är mörk,Att världen,Du perfekt harmoniOch återgå till vägen.
		-- Lao Tse, "Tao Te Ching"

%
AmbitionDe som vill förändra världenEnligt deras önskanDet går inte att lyckas.Världen formas av vägen;Det kan inte formas av jaget.Försöka förändra det, skadar du det;Försöker besittning, förlorar du den.Så några kommer att leda, medan andra följer.Vissa kommer att vara varm, andra kalltVissa kommer att vara stark, andra svaga.Vissa kommer att komma dit de skaMedan andra faller vid sidan av vägen.Så den vise blir varken extravaganta eller våldsam.
		-- Lao Tse, "Tao Te Ching"

%
VåldMäktiga män är klokt att inte använda våld,För våld har en vana att återvända;Törnen och ogräs växer överallt där en armé går,Och magra år följer ett stort krig.En allmänhet kloktFör att uppnå något mer än hans order:Inte att dra nytta av sin seger.Inte heller till ära, skryta eller stolthet själv;Att göra vad som dikteras av nödvändighet,Inte genom val.För även den starkaste kraften kommer att försvagas med tiden,Och sedan dess våld kommer att återvända, och döda den.
		-- Lao Tse, "Tao Te Ching"

%
arméerArméer är verktyg för våld;De orsakar män att hata och rädsla.Den vise kommer inte gå med dem.Hans syfte är skapelse;Deras syfte är förstörelse.Vapen är verktyg för våld,Inte av den vise;Han använder dem bara när det inte finns något val,Och sedan lugnt och med takt,För han finner ingen skönhet i dem.Den som finner skönhet i vapenDelights i slakt av män;Och som njuter i slaktDet går inte att nöja sig med fred.Så slakten måste sörjdeOch erövring firas med en begravning.
		-- Lao Tse, "Tao Te Ching"

%
formerVägen har ingen sann form,Och därför ingen kan styra det.Om en linjal kunde kontrollera vägenAllt skulle följaI samklang med sin önskan,Och söt regn skulle falla,Enkelt släckning varje törst.Vägen formas genom användning,Men då formen går förlorad.Inte hålla fast vid formerMen låt sensation flöde i världenSom en flod kurser ner till havet.
		-- Lao Tse, "Tao Te Ching"

%
förtjänsterSom förstår världen lärt;Vem förstår jaget är upplyst.Vem erövrar världen har styrka;Vem erövrar själv har harmoni;Som bestäms har syfte.Vem är nöjd har rikedom;Som försvarar sitt hem kan lång uthärda;Som överlämnar sitt hem kan överleva länge det.
		-- Lao Tse, "Tao Te Ching"

%
KontrolleraSättet flöden och ebb, skapar och förstör,Genomföra hela världen, delta i minsta detalj,Hävdar något tillbaka.Det föder allt,Även om det inte kontrollera dem;Den har inte för avsikt,Så det verkar oviktiga.Det är innehållet i allt;Även om det inte kontrollera dem;Den har inget undantag,Så det verkar ytterst viktiga.Den vise skulle inte styra världen;Han är i harmoni med världen.
		-- Lao Tse, "Tao Te Ching"

%
FredOm du erbjuder musik och matFrämlingar kan sluta med dig;Men om du är ense med vägenAlla människor i världen kommer att hålla digI säkerhet, hälsa, gemenskap och fred.Vägen saknar konst och smak;Det kan varken sett eller hört,Men dess fördelar kan inte vara uttömda.
		-- Lao Tse, "Tao Te Ching"

%
OppositionAtt minska någons inflytande, först expandera det;För att minska någons kraft, först öka den;Att störta någon, först upphöja dem;Att ta från någon, först ge dem.Detta är den finess genom vilken den svaga övervinna den starka:Fisk bör inte lämna sina djup,Och svärd bör inte lämna sina skidor.
		-- Lao Tse, "Tao Te Ching"

%
LugnVägen vidtar några åtgärder, men lämnar inget ogjort.När du acceptera dettaVärlden kommer att blomstra,I harmoni med naturen.Naturen inte har lust;Utan önskan, blir hjärtat tyst;På detta sätt hela världen görs lugn.
		-- Lao Tse, "Tao Te Ching"

%
RitualVäl etablerade hierarkier är inte lätta att rotlösa;Fåmans- övertygelser är inte lätt frigöras;Så ritual enthralls generation efter generation.Harmoni bryr sig inte om harmoni, och så naturligt uppnås;Men ritual är inriktad på harmoni, och kan därför inte uppnå den.Harmoni varken handlingar eller orsaker;Kärlek handlingar, men utan anledning;Rättvisa agerar för att tjäna anledning;Men rituella handlingar för att genomdriva anledning.När vägen försvinner, kvarstår harmoni;När harmoni försvinner, kvarstår kärlek;När kärleken är förlorad, kvarstår rättvisa;Och när rättvisa är förlorat, finns det fortfarande ritualer.Ritual är slutet av medkänsla och ärlighet,I början av förvirring;Tro är en färgstark hopp eller rädsla,I början av dårskap.Den vise går harmoni, inte genom hoppet;Han bor i frukten, inte blomman;Han accepterar substans, och ignorerar abstraktion.
		-- Lao Tse, "Tao Te Ching"

%
StödI mytiska gånger var allting helhet:Allt himlen var klar,Hela jorden var stabil,Alla bergen var fast,Alla flodbäddarna var fulla,Hela naturen var bördig,Och alla de styrande stöddes.Men att förlora klarhet, slet himlen;Förlora stabilitet, den delade jorden;Att förlora styrka, sjönk bergen;Att förlora vatten, knäckt flodbäddar;Att förlora fertilitet, försvann natur;Och förlora stöd, föll de styrande.Linjaler beroende sina undersåtar,Den ädla bero på ödmjuka;Så linjaler kallar sig föräldralösa, hungrig och ensam,För att vinna folkets stöd.
		-- Lao Tse, "Tao Te Ching"

%
Motion och användningRörelsen på vägen är att återvända;Användningen av vägen är att acceptera;Allt kommer från vägen,Och vägen kommer från ingenting.
		-- Lao Tse, "Tao Te Ching"

%
FöljandeNär den store mannen lär vägen, han följer det med flit,När den vanliga människan lär vägen, han följer det ibland;När den genomsnittliga människan lär vägen, skrattar han högt;De som inte skratta, inte lär sig alls.Därför är det sagt:Vem förstår vägen verkar dumt;Som fortskrider på vägen verkar misslyckas;Som följer vägen verkar vandra.För de finaste harmonin verkar vanligt;Den ljusaste sanning verkar färgad;Den rikaste tecken visas ofullständig;Den modigaste hjärta visas ödmjuka;Den enklaste naturen verkar obeständig.Torget, fulländade, har ingen hörn;Musik, fulländat, har ingen melodi;Kärlek, fulländade, har inget klimax;Konst, fulländat, har ingen betydelse.Vägen kan varken avkännas eller känd:Den överför sensation och överskrider kunskap.
		-- Lao Tse, "Tao Te Ching"

%
SinneVägen björnar sensation,Sensation bär minne,Sensation och minnes björn abstraktion,Och abstraktion bär hela världen;Varje sak i världen bär känsla och gör,Och genomsyras åtanke, harmoni med Way.Som andra har lärt, så gör jag undervisar,"Vem förlorar harmoni motsätter natur";Detta är roten till min undervisning.
		-- Lao Tse, "Tao Te Ching"

%
övervinnaVatten övervinner stenen;Utan ämne det kräver ingen öppning;Detta är fördelen med att vidta några åtgärder.Ändå nytta utan handling,Och erfarenhet utan abstraktion,Praktiseras av mycket få.
		-- Lao Tse, "Tao Te Ching"

%
BelåtenhetHälsa eller rykte: som hålls dyrare?Hälsa eller ägodelar: som har mer värd?Vinst eller förlust: vilket är mer besvärande?Stora kärlek medför stora kostnader,Och stor rikedom medför stor rädsla,Men belåtenhet kommer utan kostnad.För vem vet när du ska slutaFortsätter inte i fara,Och så kan länge uthärda.
		-- Lao Tse, "Tao Te Ching"

%
TystStor perfektion verkar ofullständig,Men inte förfalla;Stort överflöd verkar tom,Men inte misslyckas.Stor sanning verkar motsägelsefullt;Stor skicklighet verkar dum;Stor vältalighet verkar krångligt.När våren vinner kylan,Och hösten vinner värmen,Så lugn och tyst övervinna världen.
		-- Lao Tse, "Tao Te Ching"

%
hästarNär en nation följer vägen,Hästar bära gödsel genom sina fält;När en nation ignorerar vägen,Hästar bära soldater genom dess gator.Det finns ingen större misstag än följande önskan;Det finns ingen större katastrof än glömma belåtenhet;Det finns ingen större sjukdom än att försöka uppnå;Men en som nöjer sig med att tillfredsställa sina behovKonstaterar att belåtenhet varar.
		-- Lao Tse, "Tao Te Ching"

%
MenandeUtan att ta ett steg utomhusDu vet hela världen;Utan att ta en peep ut genom fönstretDu vet färgen på himlen.Ju mer du upplever,Ju mindre du vet.Den vise vandrar utan att veta,Ser utan att se,Åstadkommer utan att agera.
		-- Lao Tse, "Tao Te Ching"

%
OverksamhetEfterföljaren av kunskap lär så mycket som han kan varje dag;Efterföljaren på vägen glömmer så mycket som han kan varje dag.Genom avgång han når ett tillstånd av passivitetVari han gör ingenting, men ingenting återstår ogjort.Att erövra världen, uträtta någonting;Om du måste utföra något,Världen är fortfarande bortom erövring.
		-- Lao Tse, "Tao Te Ching"

%
PersonerDen vise skiljer inte mellan sig själv och världen;Behoven hos andra människor är som sin egen.Han är bra för dem som är bra;Han är också bra för dem som inte är bra,Därigenom han är bra.Han litar dem som är pålitliga;Han litar också de som inte är trovärdig,Därigenom han är pålitlig.Den vise bor i harmoni med världen,Och hans sinne är världens sinne.Så han vårdar världar andrasSom en mor gör sina barn.
		-- Lao Tse, "Tao Te Ching"

%
DödMän strömma in livet, och ebb i döden.Vissa är fyllda med livet;Vissa är tom med döden;Vissa håller fast vid livet, och därmed förgås,För livet är en abstraktion.De som är fyllda med livetBehöver inte frukta tigrar och noshörningar i vildmarken,Inte heller bära rustning och sköldar i strid;Noshörningen finner ingen plats i dem för dess horn,Tigern ingen plats för sin klo,Soldaten ingen plats för ett vapen,För döden finner ingen plats i dem.
		-- Lao Tse, "Tao Te Ching"

%
UppfostranVägen bär allt,Harmoni vårdar dem;Naturen formar dem;Användning avslutar dem.Varje följer vägen och utmärkelser harmoni,Inte enligt lag,Men genom att vara.Vägen björnar, Vårdar, former, avslutar,Skyddsrum, tröstar, och gör ett hem för dem.Bärande utan att inneha,Vårda utan tämja,Forma utan att tvinga,Detta är harmoni.
		-- Lao Tse, "Tao Te Ching"

%
KlarhetUrsprunget av världen är dess mor,Förstå mor, och du förstår barnet;Omfamna barn, och du omfamna modern,Vem kommer inte förgås när du dör.Boka dina domar och ordOch du behålla din inflytande;Säg vad du tycker och ta positionerOch ingenting kommer att spara.Som observera detalj är klarhet,Så upprätthålla flexibilitet är styrka;Använd ljuset men kasta något ljus,Så att du gör själv ingen skada,Men omfamna klarhet.
		-- Lao Tse, "Tao Te Ching"

%
svåra PathsMed men en liten förståelseMan kan följa vägen som en huvudgata,bara rädd för att lämna det;Efter en huvudgata är lätt,Ändå människor glädje i svåra banor.När palats hållsFält lämnas till ogräsOch spannmål tom;Iklädd fina kläder,Bärande vassa svärd,Glutting med mat och dryck,Hamstring rikedom och ägodelar -Dessa är de sätt för stöld,Och långt från vägen.
		-- Lao Tse, "Tao Te Ching"

%
odla HarmonyOdla harmoni inom dig själv, och harmoni blir verklig;Odla harmoni inom familjen, och harmoni blir bördig;Odla harmoni i ditt samhälle, och harmoni blirriklig;Odla harmoni i din kultur, och harmoni blirbestående;Odla harmoni i världen, och harmoni blir allestädes närvarande.Leva med en person att förstå den personen;Bo med en familj att förstå att familjen;Leva med en gemenskap för att förstå att samhället;Leva med en kultur att förstå att kulturen;Leva med världen för att förstå världen.Hur kan jag leva med världen?Genom att acceptera.
		-- Lao Tse, "Tao Te Ching"

%
mjuka BonesSom är fylld med harmoni är som en nyfödd.Getingar och ormar kommer inte bita honom;Hökar och tigrar kommer inte klo honom.Hans ben är mjuka men hans grepp är säker,För hans kött är smidig;Hans sinne är oskyldig men hans kropp är virile,För hans styrka är riklig;Hans sång är långvarig men hans röst är söt,För hans nåd är perfekt.Men att veta harmoni skapar abstraktion,Och efter abstraktion skapar ritual.Överstiger naturen skapar olycka,Och styra naturen skapar våld.
		-- Lao Tse, "Tao Te Ching"

%
OpartiskhetVem förstår inte predika;Som predikar inte förstår.Boka dina domar och ord;Släta skillnader och förlåta motsättningar;Dull din intelligens och förenkla ditt syfte;Acceptera världen.Sedan,Vänskap och fiendskap,Vinst och förlust,Ära och skam,Kommer inte att påverka dig;Världen kommer att acceptera dig.
		-- Lao Tse, "Tao Te Ching"

%
Erövra med PassivitetInte styra människor med lagar,Inte heller våld eller spioneri,Men besegra dem med passivitet.För:Ju fler moral och tabun som finns,Ju mer grymhet drabbar människor;Ju fler vapen och knivar finns,Ju fler fraktioner dela in människor;Ju fler konst och färdigheter finns,Ju mer förändring föråldrat människor;Ju fler lagar och skatter som finns,Ju mer stöld korrumperar människor.Ändå inte vidta några åtgärder, och folket vårda varandra;Gör inga lagar, och människor hanterar rättvist med varandra;Äger inget intresse, och folk samarbetar med varandra;Uttrycka ingen lust, och människorna harmonisera med varandra.
		-- Lao Tse, "Tao Te Ching"

%
No EndNär regeringen är lat och informellaMänniskorna är vänliga och ärliga;När regeringen är effektiv och svårFolket är missnöjda och bedrägliga.Turen följer på katastrof;Katastrof lurar inom lycka;Vem kan säga hur det kommer att sluta?Kanske det finns inget slut.Ärlighet är alltid lurad;Vänlighet någonsin förförd;Män har varit så här under en lång tid.Så salvia är fast men inte skära,Tillspetsade men inte piercing,Rak men inte styva,Ljusa men inte bländande.
		-- Lao Tse, "Tao Te Ching"

%
ÅterhållsamhetHantera en stor nation som du skulle laga en delikat fisk.Att styra män i enlighet med naturenDet är bäst att vara återhållsamma,Återhållsamhet gör avtal lätt att uppnå,Och lätt överenskommelse bygger harmoniska relationer;Med tillräcklig harmoni inget motstånd uppstår;När inget motstånd uppstår, då du har hjärtat avnation,Och när du har nationens hjärta, ditt inflytande kommer längehärda ut:Djupt rotad och etablerat.Detta är metoden för långt sikte och lång livslängd.
		-- Lao Tse, "Tao Te Ching"

%
demonerNär du använder vägen för att erövra världen,Dina demoner kommer att förlora sin makt för att skada.Det är inte att de förlorar sin makt som sådan,Men att de inte kommer att skada andra;Eftersom de inte kommer att skada andra,Du kommer inte att skada andra:När varken du eller dina demoner kan göra skada,Du kommer att vara i fred med dem.
		-- Lao Tse, "Tao Te Ching"

%
UnderkastelseEn nation är som en hierarki, en marknadsplats, och en jungfru.En jungfru vinner sin make genom att skicka in sina framsteg;Underkastelse är ett medel för union.Så när ett stort land underkastar sig ett litet landDet kommer att anta det lilla landet;När ett litet land underkastar sig ett stort landDet kommer att antas av det stora landet;Den lämnar och antar;De andra anfört och antas.Det är av intresse för ett stort land att förena och få service,Och i syfte att ett litet land att förena och få beskydd;Om båda skulle tjäna deras intressen,Båda måste lämna.
		-- Lao Tse, "Tao Te Ching"

%
SyndVägen är öde män,Skatten av helgonet,Och tillflykt syndaren.Fina ord är ofta lånade,Och stordåd ofta disponeras;Därför, när en man faller, inte överge honom,Och när en man vinner makt, inte hedra honom;Endast förbli opartisk och visa honom vägen.Varför skulle någon uppskattar vägen?Den gamle sade: "Genom den kan de som söker lätt att hitta,Och de som ångrar kan enkelt frikänna "Så det är den mest värdefulla gåva.
		-- Lao Tse, "Tao Te Ching"

%
SvårighetÖva ingen åtgärd;Delta göra-ingenting;Smaka på smaklös,Tora den lilla,Multiplicera fåtal,Återvända kärlek till hat.Itu med svåra medan det är ändå lätt;Ta itu med stor när det är ännu liten;Den svåra utvecklas naturligt från det enkla,Och den stora från den lilla;Så salvia, genom att behandla den lilla,Uppnår den stora.Som finner det lätt att lova har svårt att lita på;Vem tar saker lätt finner det svårt;Den vise känner igen svårigheter, och så har ingen.
		-- Lao Tse, "Tao Te Ching"

%
Skötsel i börjanVad ligger fortfarande är lätt att förstå;Vad ligger långt borta är lätt att förutse,Vad är spröd är lätt att splittras;Vad är små är lätt att sprida.Ännu ett träd bredare än en människa kan omfatta är född av en liten skott;En fördämning som är större än en flod kan svämma börjar med en klump avjord;En resa på tusen miles börjar vid plats enligt sina fötter.Därför ta itu med saker innan de inträffar;Skapa ordning innan det råder förvirring.
		-- Lao Tse, "Tao Te Ching"

%
Bryr sig slutetHan som agerar, bytet;Den som griper, förlorar.Folk misslyckas ofta på gränsen till framgång;Var försiktig i slutet som i början,Så att du kan undvika fel.Den vise önskar ingen lust,Värden no-värde,Lär ingen inlärning,Och återgår till de platser som människor har glömt;Han skulle hjälpa alla människor att bli naturligt,Men då han inte skulle vara naturlig.
		-- Lao Tse, "Tao Te Ching"

%
SubtilitetDe gamle inte försöka styra människor med kunskap,Men för att hjälpa dem att bli naturligt.Det är svårt för kunniga människor att bli naturligt.Att använda lagen för att styra en nation försvagar nationen.Men att använda naturen för att styra en nation förstärker nationen.Att förstå dessa två vägar är förståelse finess;Finess går på djupet, varierar brett,Löser förvirring och bevarar fred.
		-- Lao Tse, "Tao Te Ching"

%
Bly genom att följaFloden skär ut i dalen genom att flöda under den.Därigenom floden är herre över dalen.För att bemästra folkMan måste tala som sin tjänare;För att leda människorMan måste följa dem.Så när den vise stiger över folket,De känner sig inte förtryckta;Och när den vise står inför folket,De känner sig inte hindras.Så populariteten av salvia inte misslyckas,Han har inte påstått, och ingen har hävdat mot honom.
		-- Lao Tse, "Tao Te Ching"

%
saknar betydelseHela världen säger,"Jag är viktigt;Jag är skild från hela världen.Jag är viktigt eftersom jag är separat,Var jag samma, jag kunde aldrig vara viktigt. "Men här är tre skatterAtt jag vårda och rekommenderar till dig:Den första är medlidande,Genom vilken man finner mod.Den andra är återhållsamhet,Genom vilken en finner styrka.Och den tredje är saknar betydelse,Genom vilken man finner inflytande.De som är orädd, men utan medkänsla,Kraftfull, men utan begränsning,Eller inflytelserik, men viktigt,Det går inte att uthärda.
		-- Lao Tse, "Tao Te Ching"

%
MedlidandeMedkänsla är den finaste vapen och bästa försvaret.Om du vill skapa harmoni,Medlidande måste omge dig som en fästning.Därför,En bra soldat inger inte fruktan;En bra fighter visas inte aggression;En bra erövrare inte engagera sig i strid;En bra ledare inte utöva auktoritet.Detta är värdet av saknar betydelse;Detta är hur man vinner i samarbete med andra;Detta för hur man bygger samma harmoni som är i naturen.
		-- Lao Tse, "Tao Te Ching"

%
BakhållDet finns ett talesätt bland soldater:Det är lättare att förlora en gård än att ta en tum.På detta sätt kan man sätta in trupper utan range dem,Föra vapen för att bära utan att utsätta dem,Engagera fienden utan att invadera dem,Och uttömma sin styrka utan att bekämpa dem.Det finns ingen värre katastrof än missförstånd din fiende;För att göra detta äventyrar alla mina skatter;Så när två väl matchade krafter emot varandra,Den allmänna som underhåller medkänsla kommer att vinna.
		-- Lao Tse, "Tao Te Ching"

%
IndividualitetMina ord är lätta att förståOch mina handlingar är lätta att utföraMen ingen annan kan förstå eller utföra dem.Mina ord har betydelse; mina handlingar har anledning;Ändå dessa kan inte vara känd och jag kan inte vara känd.Vi är varje unik, och därför värdefull;Även den vise bär grova kläder, är hans hjärta jade.
		-- Lao Tse, "Tao Te Ching"

%
BegränsningSom erkänner sina begränsningar är friska,Som ignorerar sina begränsningar är sjuk.Den vise känner igen denna sjukdom som en begränsning.Och så blir immun.
		-- Lao Tse, "Tao Te Ching"

%
RotationNär folk har inget mer att förlora,Sedan revolutionen kommer att leda till.Ta inte bort sina marker,Och inte förstöra deras försörjning;Om din börda är inte tung då de inte kommer dra sig undan det.Den vise håller sig men avkräver ingen hyllning,Värden själv men kräver inga ära;Han ignorerar abstraktion och accepterar substans.
		-- Lao Tse, "Tao Te Ching"

%
ÖdeVem är modig och djärv kommer att förgås;Vem är modig och subtil kommer att gynnas.Den subtila vinst där fet förgåsFör Ödet inte hedra vågad.Och även den vise inte vågar utmana ödet.Ödet inte attackera, men alla saker erövras av det;Det är inte fråga, men alla saker svara på det;Det kallar inte, men alla saker möter den;Det är inte planera, men allt bestäms av det.Ödet netto är omfattande och mask är grov,Men ingen undkomma den.
		-- Lao Tse, "Tao Te Ching"

%
UtförandeOm människor inte rädd för döden,Vad skulle vara användningen av en bödel?Om folk bara var rädd för döden,Och du utförde alla som inte lyder,Ingen skulle våga att inte lyda dig.Vad skulle vara användningen av en bödel?Människor fruktar döden, eftersom döden är ett instrument för ödet.När människor dödas genom avrättning snarare än av ödet,Det är som carving trä i stället för en snickare.De som rista trä i stället för en snickareOfta skadar sina händer.
		-- Lao Tse, "Tao Te Ching"

%
UpprorNär linjaler ta fiberriktningen så att de kan festa,Deras människor blir hungrig;När linjaler vidta åtgärder för att tjäna sina egna intressen,Deras människor blir upprorisk;När linjaler ta liv så att deras egna liv upprätthålls,Deras människor inte längre fruktar döden.När människor agerar utan hänsyn till sina egna livDe övervinna dem som värdesätter bara sina egna liv.
		-- Lao Tse, "Tao Te Ching"

%
FlexibilitetEn nyfödd är mjuk och anbud,En crone, hård och stel.Växter och djur, i livet, är smidig och saftiga;I döden, vissnade och torr.Så mjukhet och ömhet är attribut i livet,Och hårdhet och styvhet, attribut döden.Precis som en TORR träd kommer att dela och förfallSå en oflexibel kraft kommer att möta nederlag;Den hårda och mäktig lie under markytanMedan anbud och svaga dans på vinden ovanför.
		-- Lao Tse, "Tao Te Ching"

%
BehovÄr verkan av naturen inte olikt som drar en pilbåge?Vad är högre dras ned, och vad är lägre höjs upp;Vad är högre förkortas, och vad som är tunnare breddas;Naturens rörelse minskar dem som har mer än de behöverOch ökar dem som behöver mer än de har.Det är inte så med människan.Man minskar dem som behöver mer än de harOch ökar dem som har mer än de behöver.Att ge bort vad du inte behöver är att följa vägen.Så den vise ger utan förväntan,Åstadkommer utan att kräva kredit,Och har ingen önskan om prål.
		-- Lao Tse, "Tao Te Ching"

%
vilket gavIngenting i världen är så mjuk och ger som vatten,Ändå ingenting kan bättre övervinna den hårda och starka,För de kan inte kontrollera eller göra sig av med det.Den mjuka övervinner det hårda,Den eftergivlig övervinner den starka;Varje person som känner till detta,Men ingen kan utöva den.Vem sköter folk skulle styra landet och spannmål;Vem sköter staten skulle kontrollera hela världen;Sanningen är lätt döljs av retorik.
		-- Lao Tse, "Tao Te Ching"

%
FörsoningNär konflikten stäms, några hårda känslor kvar;Detta är farligt.Den vise accepterar mindre än berorOch inte skylla eller straffa;Harmoni söker enighetDär rättvisa söker betalning.Den gamle sade: "natur är opartisk;Därför tjänar de som tjänar alla. "
		-- Lao Tse, "Tao Te Ching"

%
utopiLåt din grupp vara små, med endast ett fåtal personer,Håll verktyg i överflöd, men inte beroende av dem;Uppskattar ditt liv och vara nöjd med ditt hem;Segelbåtar och rida hästar, men inte gå för långt;Håll vapen och rustningar, men inte använda dem;Låt alla läsa och skriva,Ät gott och göra vackra saker.Leva i fred och glädje i ditt eget samhälle;Bo inom kuk-gala av dina grannar,Men behålla din självständighet från dem.
		-- Lao Tse, "Tao Te Ching"

%
The SageÄrliga människor använder ingen retorik;Retorik är inte ärlighet.Upplysta människor är inte odlas;Kultur är inte upplysning.Innehålls människor är inte rika;Rikedom är inte förnöjsamhet.Så den vise inte tjänar själv;Ju mer han gör för andra, ju mer han är nöjd;Ju mer han ger, ju mer han får.Naturen blomstrar på bekostnad av någon;Så vis gynnar alla män och har hävdat med ingen.
		-- Lao Tse, "Tao Te Ching"

%
